-- soc_system.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity soc_system is
	port (
		button_pio_external_connection_export : in    std_logic_vector(1 downto 0)  := (others => '0'); -- button_pio_external_connection.export
		clk_clk                               : in    std_logic                     := '0';             --                            clk.clk
		dipsw_pio_external_connection_export  : in    std_logic_vector(3 downto 0)  := (others => '0'); --  dipsw_pio_external_connection.export
		hps_0_h2f_reset_reset_n               : out   std_logic;                                        --                hps_0_h2f_reset.reset_n
		hps_0_hps_io_hps_io_emac1_inst_TX_CLK : out   std_logic;                                        --                   hps_0_hps_io.hps_io_emac1_inst_TX_CLK
		hps_0_hps_io_hps_io_emac1_inst_TXD0   : out   std_logic;                                        --                               .hps_io_emac1_inst_TXD0
		hps_0_hps_io_hps_io_emac1_inst_TXD1   : out   std_logic;                                        --                               .hps_io_emac1_inst_TXD1
		hps_0_hps_io_hps_io_emac1_inst_TXD2   : out   std_logic;                                        --                               .hps_io_emac1_inst_TXD2
		hps_0_hps_io_hps_io_emac1_inst_TXD3   : out   std_logic;                                        --                               .hps_io_emac1_inst_TXD3
		hps_0_hps_io_hps_io_emac1_inst_RXD0   : in    std_logic                     := '0';             --                               .hps_io_emac1_inst_RXD0
		hps_0_hps_io_hps_io_emac1_inst_MDIO   : inout std_logic                     := '0';             --                               .hps_io_emac1_inst_MDIO
		hps_0_hps_io_hps_io_emac1_inst_MDC    : out   std_logic;                                        --                               .hps_io_emac1_inst_MDC
		hps_0_hps_io_hps_io_emac1_inst_RX_CTL : in    std_logic                     := '0';             --                               .hps_io_emac1_inst_RX_CTL
		hps_0_hps_io_hps_io_emac1_inst_TX_CTL : out   std_logic;                                        --                               .hps_io_emac1_inst_TX_CTL
		hps_0_hps_io_hps_io_emac1_inst_RX_CLK : in    std_logic                     := '0';             --                               .hps_io_emac1_inst_RX_CLK
		hps_0_hps_io_hps_io_emac1_inst_RXD1   : in    std_logic                     := '0';             --                               .hps_io_emac1_inst_RXD1
		hps_0_hps_io_hps_io_emac1_inst_RXD2   : in    std_logic                     := '0';             --                               .hps_io_emac1_inst_RXD2
		hps_0_hps_io_hps_io_emac1_inst_RXD3   : in    std_logic                     := '0';             --                               .hps_io_emac1_inst_RXD3
		hps_0_hps_io_hps_io_sdio_inst_CMD     : inout std_logic                     := '0';             --                               .hps_io_sdio_inst_CMD
		hps_0_hps_io_hps_io_sdio_inst_D0      : inout std_logic                     := '0';             --                               .hps_io_sdio_inst_D0
		hps_0_hps_io_hps_io_sdio_inst_D1      : inout std_logic                     := '0';             --                               .hps_io_sdio_inst_D1
		hps_0_hps_io_hps_io_sdio_inst_CLK     : out   std_logic;                                        --                               .hps_io_sdio_inst_CLK
		hps_0_hps_io_hps_io_sdio_inst_D2      : inout std_logic                     := '0';             --                               .hps_io_sdio_inst_D2
		hps_0_hps_io_hps_io_sdio_inst_D3      : inout std_logic                     := '0';             --                               .hps_io_sdio_inst_D3
		hps_0_hps_io_hps_io_usb1_inst_D0      : inout std_logic                     := '0';             --                               .hps_io_usb1_inst_D0
		hps_0_hps_io_hps_io_usb1_inst_D1      : inout std_logic                     := '0';             --                               .hps_io_usb1_inst_D1
		hps_0_hps_io_hps_io_usb1_inst_D2      : inout std_logic                     := '0';             --                               .hps_io_usb1_inst_D2
		hps_0_hps_io_hps_io_usb1_inst_D3      : inout std_logic                     := '0';             --                               .hps_io_usb1_inst_D3
		hps_0_hps_io_hps_io_usb1_inst_D4      : inout std_logic                     := '0';             --                               .hps_io_usb1_inst_D4
		hps_0_hps_io_hps_io_usb1_inst_D5      : inout std_logic                     := '0';             --                               .hps_io_usb1_inst_D5
		hps_0_hps_io_hps_io_usb1_inst_D6      : inout std_logic                     := '0';             --                               .hps_io_usb1_inst_D6
		hps_0_hps_io_hps_io_usb1_inst_D7      : inout std_logic                     := '0';             --                               .hps_io_usb1_inst_D7
		hps_0_hps_io_hps_io_usb1_inst_CLK     : in    std_logic                     := '0';             --                               .hps_io_usb1_inst_CLK
		hps_0_hps_io_hps_io_usb1_inst_STP     : out   std_logic;                                        --                               .hps_io_usb1_inst_STP
		hps_0_hps_io_hps_io_usb1_inst_DIR     : in    std_logic                     := '0';             --                               .hps_io_usb1_inst_DIR
		hps_0_hps_io_hps_io_usb1_inst_NXT     : in    std_logic                     := '0';             --                               .hps_io_usb1_inst_NXT
		hps_0_hps_io_hps_io_spim1_inst_CLK    : out   std_logic;                                        --                               .hps_io_spim1_inst_CLK
		hps_0_hps_io_hps_io_spim1_inst_MOSI   : out   std_logic;                                        --                               .hps_io_spim1_inst_MOSI
		hps_0_hps_io_hps_io_spim1_inst_MISO   : in    std_logic                     := '0';             --                               .hps_io_spim1_inst_MISO
		hps_0_hps_io_hps_io_spim1_inst_SS0    : out   std_logic;                                        --                               .hps_io_spim1_inst_SS0
		hps_0_hps_io_hps_io_uart0_inst_RX     : in    std_logic                     := '0';             --                               .hps_io_uart0_inst_RX
		hps_0_hps_io_hps_io_uart0_inst_TX     : out   std_logic;                                        --                               .hps_io_uart0_inst_TX
		hps_0_hps_io_hps_io_i2c0_inst_SDA     : inout std_logic                     := '0';             --                               .hps_io_i2c0_inst_SDA
		hps_0_hps_io_hps_io_i2c0_inst_SCL     : inout std_logic                     := '0';             --                               .hps_io_i2c0_inst_SCL
		hps_0_hps_io_hps_io_i2c1_inst_SDA     : inout std_logic                     := '0';             --                               .hps_io_i2c1_inst_SDA
		hps_0_hps_io_hps_io_i2c1_inst_SCL     : inout std_logic                     := '0';             --                               .hps_io_i2c1_inst_SCL
		hps_0_hps_io_hps_io_gpio_inst_GPIO09  : inout std_logic                     := '0';             --                               .hps_io_gpio_inst_GPIO09
		hps_0_hps_io_hps_io_gpio_inst_GPIO35  : inout std_logic                     := '0';             --                               .hps_io_gpio_inst_GPIO35
		hps_0_hps_io_hps_io_gpio_inst_GPIO40  : inout std_logic                     := '0';             --                               .hps_io_gpio_inst_GPIO40
		hps_0_hps_io_hps_io_gpio_inst_GPIO53  : inout std_logic                     := '0';             --                               .hps_io_gpio_inst_GPIO53
		hps_0_hps_io_hps_io_gpio_inst_GPIO54  : inout std_logic                     := '0';             --                               .hps_io_gpio_inst_GPIO54
		hps_0_hps_io_hps_io_gpio_inst_GPIO61  : inout std_logic                     := '0';             --                               .hps_io_gpio_inst_GPIO61
		ip_servomotor_0_conduit_end_commande  : out   std_logic;                                        --    ip_servomotor_0_conduit_end.commande
		ip_servomotor_0_conduit_end_led       : out   std_logic_vector(7 downto 0);                     --                               .led
		led_pio_external_connection_export    : out   std_logic_vector(7 downto 0);                     --    led_pio_external_connection.export
		memory_mem_a                          : out   std_logic_vector(14 downto 0);                    --                         memory.mem_a
		memory_mem_ba                         : out   std_logic_vector(2 downto 0);                     --                               .mem_ba
		memory_mem_ck                         : out   std_logic;                                        --                               .mem_ck
		memory_mem_ck_n                       : out   std_logic;                                        --                               .mem_ck_n
		memory_mem_cke                        : out   std_logic;                                        --                               .mem_cke
		memory_mem_cs_n                       : out   std_logic;                                        --                               .mem_cs_n
		memory_mem_ras_n                      : out   std_logic;                                        --                               .mem_ras_n
		memory_mem_cas_n                      : out   std_logic;                                        --                               .mem_cas_n
		memory_mem_we_n                       : out   std_logic;                                        --                               .mem_we_n
		memory_mem_reset_n                    : out   std_logic;                                        --                               .mem_reset_n
		memory_mem_dq                         : inout std_logic_vector(31 downto 0) := (others => '0'); --                               .mem_dq
		memory_mem_dqs                        : inout std_logic_vector(3 downto 0)  := (others => '0'); --                               .mem_dqs
		memory_mem_dqs_n                      : inout std_logic_vector(3 downto 0)  := (others => '0'); --                               .mem_dqs_n
		memory_mem_odt                        : out   std_logic;                                        --                               .mem_odt
		memory_mem_dm                         : out   std_logic_vector(3 downto 0);                     --                               .mem_dm
		memory_oct_rzqin                      : in    std_logic                     := '0';             --                               .oct_rzqin
		reset_reset_n                         : in    std_logic                     := '0'              --                          reset.reset_n
	);
end entity soc_system;

architecture rtl of soc_system is
	component DF9GMS is
		generic (
			Fclock : positive := 50000000
		);
		port (
			address     : in  std_logic                    := 'X';             -- address
			write_data  : in  std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			write_n     : in  std_logic                    := 'X';             -- write_n
			chip_select : in  std_logic                    := 'X';             -- chipselect
			CLK         : in  std_logic                    := 'X';             -- clk
			pulse       : out std_logic;                                       -- commande
			led         : out std_logic_vector(7 downto 0);                    -- led
			RST_n       : in  std_logic                    := 'X'              -- reset_n
		);
	end component DF9GMS;

	component soc_system_button_pio is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component soc_system_button_pio;

	component soc_system_d is
		generic (
			F2S_Width : integer := 2;
			S2F_Width : integer := 2
		);
		port (
			mem_a                    : out   std_logic_vector(14 downto 0);                     -- mem_a
			mem_ba                   : out   std_logic_vector(2 downto 0);                      -- mem_ba
			mem_ck                   : out   std_logic;                                         -- mem_ck
			mem_ck_n                 : out   std_logic;                                         -- mem_ck_n
			mem_cke                  : out   std_logic;                                         -- mem_cke
			mem_cs_n                 : out   std_logic;                                         -- mem_cs_n
			mem_ras_n                : out   std_logic;                                         -- mem_ras_n
			mem_cas_n                : out   std_logic;                                         -- mem_cas_n
			mem_we_n                 : out   std_logic;                                         -- mem_we_n
			mem_reset_n              : out   std_logic;                                         -- mem_reset_n
			mem_dq                   : inout std_logic_vector(31 downto 0)  := (others => 'X'); -- mem_dq
			mem_dqs                  : inout std_logic_vector(3 downto 0)   := (others => 'X'); -- mem_dqs
			mem_dqs_n                : inout std_logic_vector(3 downto 0)   := (others => 'X'); -- mem_dqs_n
			mem_odt                  : out   std_logic;                                         -- mem_odt
			mem_dm                   : out   std_logic_vector(3 downto 0);                      -- mem_dm
			oct_rzqin                : in    std_logic                      := 'X';             -- oct_rzqin
			hps_io_emac1_inst_TX_CLK : out   std_logic;                                         -- hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   : out   std_logic;                                         -- hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   : out   std_logic;                                         -- hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   : out   std_logic;                                         -- hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   : out   std_logic;                                         -- hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   : inout std_logic                      := 'X';             -- hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    : out   std_logic;                                         -- hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL : out   std_logic;                                         -- hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RXD3
			hps_io_sdio_inst_CMD     : inout std_logic                      := 'X';             -- hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      : inout std_logic                      := 'X';             -- hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      : inout std_logic                      := 'X';             -- hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     : out   std_logic;                                         -- hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      : inout std_logic                      := 'X';             -- hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      : inout std_logic                      := 'X';             -- hps_io_sdio_inst_D3
			hps_io_usb1_inst_D0      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D0
			hps_io_usb1_inst_D1      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D1
			hps_io_usb1_inst_D2      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D2
			hps_io_usb1_inst_D3      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D3
			hps_io_usb1_inst_D4      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D4
			hps_io_usb1_inst_D5      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D5
			hps_io_usb1_inst_D6      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D6
			hps_io_usb1_inst_D7      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D7
			hps_io_usb1_inst_CLK     : in    std_logic                      := 'X';             -- hps_io_usb1_inst_CLK
			hps_io_usb1_inst_STP     : out   std_logic;                                         -- hps_io_usb1_inst_STP
			hps_io_usb1_inst_DIR     : in    std_logic                      := 'X';             -- hps_io_usb1_inst_DIR
			hps_io_usb1_inst_NXT     : in    std_logic                      := 'X';             -- hps_io_usb1_inst_NXT
			hps_io_spim1_inst_CLK    : out   std_logic;                                         -- hps_io_spim1_inst_CLK
			hps_io_spim1_inst_MOSI   : out   std_logic;                                         -- hps_io_spim1_inst_MOSI
			hps_io_spim1_inst_MISO   : in    std_logic                      := 'X';             -- hps_io_spim1_inst_MISO
			hps_io_spim1_inst_SS0    : out   std_logic;                                         -- hps_io_spim1_inst_SS0
			hps_io_uart0_inst_RX     : in    std_logic                      := 'X';             -- hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     : out   std_logic;                                         -- hps_io_uart0_inst_TX
			hps_io_i2c0_inst_SDA     : inout std_logic                      := 'X';             -- hps_io_i2c0_inst_SDA
			hps_io_i2c0_inst_SCL     : inout std_logic                      := 'X';             -- hps_io_i2c0_inst_SCL
			hps_io_i2c1_inst_SDA     : inout std_logic                      := 'X';             -- hps_io_i2c1_inst_SDA
			hps_io_i2c1_inst_SCL     : inout std_logic                      := 'X';             -- hps_io_i2c1_inst_SCL
			hps_io_gpio_inst_GPIO09  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO09
			hps_io_gpio_inst_GPIO35  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO35
			hps_io_gpio_inst_GPIO40  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO40
			hps_io_gpio_inst_GPIO53  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO53
			hps_io_gpio_inst_GPIO54  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO54
			hps_io_gpio_inst_GPIO61  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO61
			h2f_rst_n                : out   std_logic;                                         -- reset_n
			h2f_axi_clk              : in    std_logic                      := 'X';             -- clk
			h2f_AWID                 : out   std_logic_vector(11 downto 0);                     -- awid
			h2f_AWADDR               : out   std_logic_vector(29 downto 0);                     -- awaddr
			h2f_AWLEN                : out   std_logic_vector(3 downto 0);                      -- awlen
			h2f_AWSIZE               : out   std_logic_vector(2 downto 0);                      -- awsize
			h2f_AWBURST              : out   std_logic_vector(1 downto 0);                      -- awburst
			h2f_AWLOCK               : out   std_logic_vector(1 downto 0);                      -- awlock
			h2f_AWCACHE              : out   std_logic_vector(3 downto 0);                      -- awcache
			h2f_AWPROT               : out   std_logic_vector(2 downto 0);                      -- awprot
			h2f_AWVALID              : out   std_logic;                                         -- awvalid
			h2f_AWREADY              : in    std_logic                      := 'X';             -- awready
			h2f_WID                  : out   std_logic_vector(11 downto 0);                     -- wid
			h2f_WDATA                : out   std_logic_vector(63 downto 0);                     -- wdata
			h2f_WSTRB                : out   std_logic_vector(7 downto 0);                      -- wstrb
			h2f_WLAST                : out   std_logic;                                         -- wlast
			h2f_WVALID               : out   std_logic;                                         -- wvalid
			h2f_WREADY               : in    std_logic                      := 'X';             -- wready
			h2f_BID                  : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- bid
			h2f_BRESP                : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- bresp
			h2f_BVALID               : in    std_logic                      := 'X';             -- bvalid
			h2f_BREADY               : out   std_logic;                                         -- bready
			h2f_ARID                 : out   std_logic_vector(11 downto 0);                     -- arid
			h2f_ARADDR               : out   std_logic_vector(29 downto 0);                     -- araddr
			h2f_ARLEN                : out   std_logic_vector(3 downto 0);                      -- arlen
			h2f_ARSIZE               : out   std_logic_vector(2 downto 0);                      -- arsize
			h2f_ARBURST              : out   std_logic_vector(1 downto 0);                      -- arburst
			h2f_ARLOCK               : out   std_logic_vector(1 downto 0);                      -- arlock
			h2f_ARCACHE              : out   std_logic_vector(3 downto 0);                      -- arcache
			h2f_ARPROT               : out   std_logic_vector(2 downto 0);                      -- arprot
			h2f_ARVALID              : out   std_logic;                                         -- arvalid
			h2f_ARREADY              : in    std_logic                      := 'X';             -- arready
			h2f_RID                  : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- rid
			h2f_RDATA                : in    std_logic_vector(63 downto 0)  := (others => 'X'); -- rdata
			h2f_RRESP                : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- rresp
			h2f_RLAST                : in    std_logic                      := 'X';             -- rlast
			h2f_RVALID               : in    std_logic                      := 'X';             -- rvalid
			h2f_RREADY               : out   std_logic;                                         -- rready
			f2h_axi_clk              : in    std_logic                      := 'X';             -- clk
			f2h_AWID                 : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- awid
			f2h_AWADDR               : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- awaddr
			f2h_AWLEN                : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- awlen
			f2h_AWSIZE               : in    std_logic_vector(2 downto 0)   := (others => 'X'); -- awsize
			f2h_AWBURST              : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- awburst
			f2h_AWLOCK               : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- awlock
			f2h_AWCACHE              : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- awcache
			f2h_AWPROT               : in    std_logic_vector(2 downto 0)   := (others => 'X'); -- awprot
			f2h_AWVALID              : in    std_logic                      := 'X';             -- awvalid
			f2h_AWREADY              : out   std_logic;                                         -- awready
			f2h_AWUSER               : in    std_logic_vector(4 downto 0)   := (others => 'X'); -- awuser
			f2h_WID                  : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- wid
			f2h_WDATA                : in    std_logic_vector(127 downto 0) := (others => 'X'); -- wdata
			f2h_WSTRB                : in    std_logic_vector(15 downto 0)  := (others => 'X'); -- wstrb
			f2h_WLAST                : in    std_logic                      := 'X';             -- wlast
			f2h_WVALID               : in    std_logic                      := 'X';             -- wvalid
			f2h_WREADY               : out   std_logic;                                         -- wready
			f2h_BID                  : out   std_logic_vector(7 downto 0);                      -- bid
			f2h_BRESP                : out   std_logic_vector(1 downto 0);                      -- bresp
			f2h_BVALID               : out   std_logic;                                         -- bvalid
			f2h_BREADY               : in    std_logic                      := 'X';             -- bready
			f2h_ARID                 : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- arid
			f2h_ARADDR               : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- araddr
			f2h_ARLEN                : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- arlen
			f2h_ARSIZE               : in    std_logic_vector(2 downto 0)   := (others => 'X'); -- arsize
			f2h_ARBURST              : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- arburst
			f2h_ARLOCK               : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- arlock
			f2h_ARCACHE              : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- arcache
			f2h_ARPROT               : in    std_logic_vector(2 downto 0)   := (others => 'X'); -- arprot
			f2h_ARVALID              : in    std_logic                      := 'X';             -- arvalid
			f2h_ARREADY              : out   std_logic;                                         -- arready
			f2h_ARUSER               : in    std_logic_vector(4 downto 0)   := (others => 'X'); -- aruser
			f2h_RID                  : out   std_logic_vector(7 downto 0);                      -- rid
			f2h_RDATA                : out   std_logic_vector(127 downto 0);                    -- rdata
			f2h_RRESP                : out   std_logic_vector(1 downto 0);                      -- rresp
			f2h_RLAST                : out   std_logic;                                         -- rlast
			f2h_RVALID               : out   std_logic;                                         -- rvalid
			f2h_RREADY               : in    std_logic                      := 'X';             -- rready
			h2f_lw_axi_clk           : in    std_logic                      := 'X';             -- clk
			h2f_lw_AWID              : out   std_logic_vector(11 downto 0);                     -- awid
			h2f_lw_AWADDR            : out   std_logic_vector(20 downto 0);                     -- awaddr
			h2f_lw_AWLEN             : out   std_logic_vector(3 downto 0);                      -- awlen
			h2f_lw_AWSIZE            : out   std_logic_vector(2 downto 0);                      -- awsize
			h2f_lw_AWBURST           : out   std_logic_vector(1 downto 0);                      -- awburst
			h2f_lw_AWLOCK            : out   std_logic_vector(1 downto 0);                      -- awlock
			h2f_lw_AWCACHE           : out   std_logic_vector(3 downto 0);                      -- awcache
			h2f_lw_AWPROT            : out   std_logic_vector(2 downto 0);                      -- awprot
			h2f_lw_AWVALID           : out   std_logic;                                         -- awvalid
			h2f_lw_AWREADY           : in    std_logic                      := 'X';             -- awready
			h2f_lw_WID               : out   std_logic_vector(11 downto 0);                     -- wid
			h2f_lw_WDATA             : out   std_logic_vector(31 downto 0);                     -- wdata
			h2f_lw_WSTRB             : out   std_logic_vector(3 downto 0);                      -- wstrb
			h2f_lw_WLAST             : out   std_logic;                                         -- wlast
			h2f_lw_WVALID            : out   std_logic;                                         -- wvalid
			h2f_lw_WREADY            : in    std_logic                      := 'X';             -- wready
			h2f_lw_BID               : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- bid
			h2f_lw_BRESP             : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- bresp
			h2f_lw_BVALID            : in    std_logic                      := 'X';             -- bvalid
			h2f_lw_BREADY            : out   std_logic;                                         -- bready
			h2f_lw_ARID              : out   std_logic_vector(11 downto 0);                     -- arid
			h2f_lw_ARADDR            : out   std_logic_vector(20 downto 0);                     -- araddr
			h2f_lw_ARLEN             : out   std_logic_vector(3 downto 0);                      -- arlen
			h2f_lw_ARSIZE            : out   std_logic_vector(2 downto 0);                      -- arsize
			h2f_lw_ARBURST           : out   std_logic_vector(1 downto 0);                      -- arburst
			h2f_lw_ARLOCK            : out   std_logic_vector(1 downto 0);                      -- arlock
			h2f_lw_ARCACHE           : out   std_logic_vector(3 downto 0);                      -- arcache
			h2f_lw_ARPROT            : out   std_logic_vector(2 downto 0);                      -- arprot
			h2f_lw_ARVALID           : out   std_logic;                                         -- arvalid
			h2f_lw_ARREADY           : in    std_logic                      := 'X';             -- arready
			h2f_lw_RID               : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- rid
			h2f_lw_RDATA             : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- rdata
			h2f_lw_RRESP             : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- rresp
			h2f_lw_RLAST             : in    std_logic                      := 'X';             -- rlast
			h2f_lw_RVALID            : in    std_logic                      := 'X';             -- rvalid
			h2f_lw_RREADY            : out   std_logic;                                         -- rready
			f2h_irq_p0               : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- irq
			f2h_irq_p1               : in    std_logic_vector(31 downto 0)  := (others => 'X')  -- irq
		);
	end component soc_system_d;

	component soc_system_dipsw_pio is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component soc_system_dipsw_pio;

	component soc_system_fpga_only_master is
		generic (
			USE_PLI     : integer := 0;
			PLI_PORT    : integer := 50000;
			FIFO_DEPTHS : integer := 2
		);
		port (
			clk_clk              : in  std_logic                     := 'X';             -- clk
			clk_reset_reset      : in  std_logic                     := 'X';             -- reset
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			master_read          : out std_logic;                                        -- read
			master_write         : out std_logic;                                        -- write
			master_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			master_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			master_reset_reset   : out std_logic                                         -- reset
		);
	end component soc_system_fpga_only_master;

	component intr_capturer is
		generic (
			NUM_INTR : integer := 32
		);
		port (
			clk          : in  std_logic                     := 'X';             -- clk
			rst_n        : in  std_logic                     := 'X';             -- reset_n
			addr         : in  std_logic                     := 'X';             -- address
			read         : in  std_logic                     := 'X';             -- read
			rddata       : out std_logic_vector(31 downto 0);                    -- readdata
			interrupt_in : in  std_logic_vector(31 downto 0) := (others => 'X')  -- irq
		);
	end component intr_capturer;

	component soc_system_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component soc_system_jtag_uart;

	component soc_system_led_pio is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component soc_system_led_pio;

	component soc_system_onchip_memory2_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(63 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(63 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component soc_system_onchip_memory2_0;

	component soc_system_sysid_qsys is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component soc_system_sysid_qsys;

	component soc_system_mm_interconnect_0 is
		port (
			d_h2f_axi_master_awid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- awid
			d_h2f_axi_master_awaddr                                      : in  std_logic_vector(29 downto 0) := (others => 'X'); -- awaddr
			d_h2f_axi_master_awlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awlen
			d_h2f_axi_master_awsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			d_h2f_axi_master_awburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			d_h2f_axi_master_awlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awlock
			d_h2f_axi_master_awcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			d_h2f_axi_master_awprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			d_h2f_axi_master_awvalid                                     : in  std_logic                     := 'X';             -- awvalid
			d_h2f_axi_master_awready                                     : out std_logic;                                        -- awready
			d_h2f_axi_master_wid                                         : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wid
			d_h2f_axi_master_wdata                                       : in  std_logic_vector(63 downto 0) := (others => 'X'); -- wdata
			d_h2f_axi_master_wstrb                                       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wstrb
			d_h2f_axi_master_wlast                                       : in  std_logic                     := 'X';             -- wlast
			d_h2f_axi_master_wvalid                                      : in  std_logic                     := 'X';             -- wvalid
			d_h2f_axi_master_wready                                      : out std_logic;                                        -- wready
			d_h2f_axi_master_bid                                         : out std_logic_vector(11 downto 0);                    -- bid
			d_h2f_axi_master_bresp                                       : out std_logic_vector(1 downto 0);                     -- bresp
			d_h2f_axi_master_bvalid                                      : out std_logic;                                        -- bvalid
			d_h2f_axi_master_bready                                      : in  std_logic                     := 'X';             -- bready
			d_h2f_axi_master_arid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- arid
			d_h2f_axi_master_araddr                                      : in  std_logic_vector(29 downto 0) := (others => 'X'); -- araddr
			d_h2f_axi_master_arlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arlen
			d_h2f_axi_master_arsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			d_h2f_axi_master_arburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			d_h2f_axi_master_arlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arlock
			d_h2f_axi_master_arcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			d_h2f_axi_master_arprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			d_h2f_axi_master_arvalid                                     : in  std_logic                     := 'X';             -- arvalid
			d_h2f_axi_master_arready                                     : out std_logic;                                        -- arready
			d_h2f_axi_master_rid                                         : out std_logic_vector(11 downto 0);                    -- rid
			d_h2f_axi_master_rdata                                       : out std_logic_vector(63 downto 0);                    -- rdata
			d_h2f_axi_master_rresp                                       : out std_logic_vector(1 downto 0);                     -- rresp
			d_h2f_axi_master_rlast                                       : out std_logic;                                        -- rlast
			d_h2f_axi_master_rvalid                                      : out std_logic;                                        -- rvalid
			d_h2f_axi_master_rready                                      : in  std_logic                     := 'X';             -- rready
			d_h2f_lw_axi_master_awid                                     : in  std_logic_vector(11 downto 0) := (others => 'X'); -- awid
			d_h2f_lw_axi_master_awaddr                                   : in  std_logic_vector(20 downto 0) := (others => 'X'); -- awaddr
			d_h2f_lw_axi_master_awlen                                    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awlen
			d_h2f_lw_axi_master_awsize                                   : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			d_h2f_lw_axi_master_awburst                                  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			d_h2f_lw_axi_master_awlock                                   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awlock
			d_h2f_lw_axi_master_awcache                                  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			d_h2f_lw_axi_master_awprot                                   : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			d_h2f_lw_axi_master_awvalid                                  : in  std_logic                     := 'X';             -- awvalid
			d_h2f_lw_axi_master_awready                                  : out std_logic;                                        -- awready
			d_h2f_lw_axi_master_wid                                      : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wid
			d_h2f_lw_axi_master_wdata                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wdata
			d_h2f_lw_axi_master_wstrb                                    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- wstrb
			d_h2f_lw_axi_master_wlast                                    : in  std_logic                     := 'X';             -- wlast
			d_h2f_lw_axi_master_wvalid                                   : in  std_logic                     := 'X';             -- wvalid
			d_h2f_lw_axi_master_wready                                   : out std_logic;                                        -- wready
			d_h2f_lw_axi_master_bid                                      : out std_logic_vector(11 downto 0);                    -- bid
			d_h2f_lw_axi_master_bresp                                    : out std_logic_vector(1 downto 0);                     -- bresp
			d_h2f_lw_axi_master_bvalid                                   : out std_logic;                                        -- bvalid
			d_h2f_lw_axi_master_bready                                   : in  std_logic                     := 'X';             -- bready
			d_h2f_lw_axi_master_arid                                     : in  std_logic_vector(11 downto 0) := (others => 'X'); -- arid
			d_h2f_lw_axi_master_araddr                                   : in  std_logic_vector(20 downto 0) := (others => 'X'); -- araddr
			d_h2f_lw_axi_master_arlen                                    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arlen
			d_h2f_lw_axi_master_arsize                                   : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			d_h2f_lw_axi_master_arburst                                  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			d_h2f_lw_axi_master_arlock                                   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arlock
			d_h2f_lw_axi_master_arcache                                  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			d_h2f_lw_axi_master_arprot                                   : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			d_h2f_lw_axi_master_arvalid                                  : in  std_logic                     := 'X';             -- arvalid
			d_h2f_lw_axi_master_arready                                  : out std_logic;                                        -- arready
			d_h2f_lw_axi_master_rid                                      : out std_logic_vector(11 downto 0);                    -- rid
			d_h2f_lw_axi_master_rdata                                    : out std_logic_vector(31 downto 0);                    -- rdata
			d_h2f_lw_axi_master_rresp                                    : out std_logic_vector(1 downto 0);                     -- rresp
			d_h2f_lw_axi_master_rlast                                    : out std_logic;                                        -- rlast
			d_h2f_lw_axi_master_rvalid                                   : out std_logic;                                        -- rvalid
			d_h2f_lw_axi_master_rready                                   : in  std_logic                     := 'X';             -- rready
			clk_0_clk_clk                                                : in  std_logic                     := 'X';             -- clk
			d_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			fpga_only_master_clk_reset_reset_bridge_in_reset_reset       : in  std_logic                     := 'X';             -- reset
			onchip_memory2_0_reset1_reset_bridge_in_reset_reset          : in  std_logic                     := 'X';             -- reset
			fpga_only_master_master_address                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			fpga_only_master_master_waitrequest                          : out std_logic;                                        -- waitrequest
			fpga_only_master_master_byteenable                           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			fpga_only_master_master_read                                 : in  std_logic                     := 'X';             -- read
			fpga_only_master_master_readdata                             : out std_logic_vector(31 downto 0);                    -- readdata
			fpga_only_master_master_readdatavalid                        : out std_logic;                                        -- readdatavalid
			fpga_only_master_master_write                                : in  std_logic                     := 'X';             -- write
			fpga_only_master_master_writedata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			button_pio_s1_address                                        : out std_logic_vector(1 downto 0);                     -- address
			button_pio_s1_write                                          : out std_logic;                                        -- write
			button_pio_s1_readdata                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			button_pio_s1_writedata                                      : out std_logic_vector(31 downto 0);                    -- writedata
			button_pio_s1_chipselect                                     : out std_logic;                                        -- chipselect
			dipsw_pio_s1_address                                         : out std_logic_vector(1 downto 0);                     -- address
			dipsw_pio_s1_write                                           : out std_logic;                                        -- write
			dipsw_pio_s1_readdata                                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			dipsw_pio_s1_writedata                                       : out std_logic_vector(31 downto 0);                    -- writedata
			dipsw_pio_s1_chipselect                                      : out std_logic;                                        -- chipselect
			intr_capturer_0_avalon_slave_0_address                       : out std_logic_vector(0 downto 0);                     -- address
			intr_capturer_0_avalon_slave_0_read                          : out std_logic;                                        -- read
			intr_capturer_0_avalon_slave_0_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			IP_Servomotor_0_avalon_slave_0_address                       : out std_logic_vector(0 downto 0);                     -- address
			IP_Servomotor_0_avalon_slave_0_write                         : out std_logic;                                        -- write
			IP_Servomotor_0_avalon_slave_0_writedata                     : out std_logic_vector(7 downto 0);                     -- writedata
			IP_Servomotor_0_avalon_slave_0_chipselect                    : out std_logic;                                        -- chipselect
			jtag_uart_avalon_jtag_slave_address                          : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write                            : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read                             : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest                      : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                       : out std_logic;                                        -- chipselect
			led_pio_s1_address                                           : out std_logic_vector(1 downto 0);                     -- address
			led_pio_s1_write                                             : out std_logic;                                        -- write
			led_pio_s1_readdata                                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			led_pio_s1_writedata                                         : out std_logic_vector(31 downto 0);                    -- writedata
			led_pio_s1_chipselect                                        : out std_logic;                                        -- chipselect
			onchip_memory2_0_s1_address                                  : out std_logic_vector(12 downto 0);                    -- address
			onchip_memory2_0_s1_write                                    : out std_logic;                                        -- write
			onchip_memory2_0_s1_readdata                                 : in  std_logic_vector(63 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_0_s1_writedata                                : out std_logic_vector(63 downto 0);                    -- writedata
			onchip_memory2_0_s1_byteenable                               : out std_logic_vector(7 downto 0);                     -- byteenable
			onchip_memory2_0_s1_chipselect                               : out std_logic;                                        -- chipselect
			onchip_memory2_0_s1_clken                                    : out std_logic;                                        -- clken
			sysid_qsys_control_slave_address                             : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_control_slave_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component soc_system_mm_interconnect_0;

	component soc_system_mm_interconnect_1 is
		port (
			d_f2h_axi_slave_awid                                                : out std_logic_vector(7 downto 0);                      -- awid
			d_f2h_axi_slave_awaddr                                              : out std_logic_vector(31 downto 0);                     -- awaddr
			d_f2h_axi_slave_awlen                                               : out std_logic_vector(3 downto 0);                      -- awlen
			d_f2h_axi_slave_awsize                                              : out std_logic_vector(2 downto 0);                      -- awsize
			d_f2h_axi_slave_awburst                                             : out std_logic_vector(1 downto 0);                      -- awburst
			d_f2h_axi_slave_awlock                                              : out std_logic_vector(1 downto 0);                      -- awlock
			d_f2h_axi_slave_awcache                                             : out std_logic_vector(3 downto 0);                      -- awcache
			d_f2h_axi_slave_awprot                                              : out std_logic_vector(2 downto 0);                      -- awprot
			d_f2h_axi_slave_awuser                                              : out std_logic_vector(4 downto 0);                      -- awuser
			d_f2h_axi_slave_awvalid                                             : out std_logic;                                         -- awvalid
			d_f2h_axi_slave_awready                                             : in  std_logic                      := 'X';             -- awready
			d_f2h_axi_slave_wid                                                 : out std_logic_vector(7 downto 0);                      -- wid
			d_f2h_axi_slave_wdata                                               : out std_logic_vector(127 downto 0);                    -- wdata
			d_f2h_axi_slave_wstrb                                               : out std_logic_vector(15 downto 0);                     -- wstrb
			d_f2h_axi_slave_wlast                                               : out std_logic;                                         -- wlast
			d_f2h_axi_slave_wvalid                                              : out std_logic;                                         -- wvalid
			d_f2h_axi_slave_wready                                              : in  std_logic                      := 'X';             -- wready
			d_f2h_axi_slave_bid                                                 : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- bid
			d_f2h_axi_slave_bresp                                               : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- bresp
			d_f2h_axi_slave_bvalid                                              : in  std_logic                      := 'X';             -- bvalid
			d_f2h_axi_slave_bready                                              : out std_logic;                                         -- bready
			d_f2h_axi_slave_arid                                                : out std_logic_vector(7 downto 0);                      -- arid
			d_f2h_axi_slave_araddr                                              : out std_logic_vector(31 downto 0);                     -- araddr
			d_f2h_axi_slave_arlen                                               : out std_logic_vector(3 downto 0);                      -- arlen
			d_f2h_axi_slave_arsize                                              : out std_logic_vector(2 downto 0);                      -- arsize
			d_f2h_axi_slave_arburst                                             : out std_logic_vector(1 downto 0);                      -- arburst
			d_f2h_axi_slave_arlock                                              : out std_logic_vector(1 downto 0);                      -- arlock
			d_f2h_axi_slave_arcache                                             : out std_logic_vector(3 downto 0);                      -- arcache
			d_f2h_axi_slave_arprot                                              : out std_logic_vector(2 downto 0);                      -- arprot
			d_f2h_axi_slave_aruser                                              : out std_logic_vector(4 downto 0);                      -- aruser
			d_f2h_axi_slave_arvalid                                             : out std_logic;                                         -- arvalid
			d_f2h_axi_slave_arready                                             : in  std_logic                      := 'X';             -- arready
			d_f2h_axi_slave_rid                                                 : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- rid
			d_f2h_axi_slave_rdata                                               : in  std_logic_vector(127 downto 0) := (others => 'X'); -- rdata
			d_f2h_axi_slave_rresp                                               : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- rresp
			d_f2h_axi_slave_rlast                                               : in  std_logic                      := 'X';             -- rlast
			d_f2h_axi_slave_rvalid                                              : in  std_logic                      := 'X';             -- rvalid
			d_f2h_axi_slave_rready                                              : out std_logic;                                         -- rready
			clk_0_clk_clk                                                       : in  std_logic                      := 'X';             -- clk
			d_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset        : in  std_logic                      := 'X';             -- reset
			hps_only_master_clk_reset_reset_bridge_in_reset_reset               : in  std_logic                      := 'X';             -- reset
			hps_only_master_master_translator_reset_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			hps_only_master_master_address                                      : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			hps_only_master_master_waitrequest                                  : out std_logic;                                         -- waitrequest
			hps_only_master_master_byteenable                                   : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			hps_only_master_master_read                                         : in  std_logic                      := 'X';             -- read
			hps_only_master_master_readdata                                     : out std_logic_vector(31 downto 0);                     -- readdata
			hps_only_master_master_readdatavalid                                : out std_logic;                                         -- readdatavalid
			hps_only_master_master_write                                        : in  std_logic                      := 'X';             -- write
			hps_only_master_master_writedata                                    : in  std_logic_vector(31 downto 0)  := (others => 'X')  -- writedata
		);
	end component soc_system_mm_interconnect_1;

	component soc_system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component soc_system_irq_mapper;

	component soc_system_irq_mapper_001 is
		port (
			clk        : in  std_logic                     := 'X'; -- clk
			reset      : in  std_logic                     := 'X'; -- reset
			sender_irq : out std_logic_vector(31 downto 0)         -- irq
		);
	end component soc_system_irq_mapper_001;

	component soc_system_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component soc_system_rst_controller;

	component soc_system_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component soc_system_rst_controller_001;

	signal d_h2f_reset_reset                                                : std_logic;                      -- d:h2f_rst_n -> [hps_0_h2f_reset_reset_n, hps_0_h2f_reset_reset_n:in]
	signal d_h2f_axi_master_awburst                                         : std_logic_vector(1 downto 0);   -- d:h2f_AWBURST -> mm_interconnect_0:d_h2f_axi_master_awburst
	signal d_h2f_axi_master_arlen                                           : std_logic_vector(3 downto 0);   -- d:h2f_ARLEN -> mm_interconnect_0:d_h2f_axi_master_arlen
	signal d_h2f_axi_master_wstrb                                           : std_logic_vector(7 downto 0);   -- d:h2f_WSTRB -> mm_interconnect_0:d_h2f_axi_master_wstrb
	signal d_h2f_axi_master_wready                                          : std_logic;                      -- mm_interconnect_0:d_h2f_axi_master_wready -> d:h2f_WREADY
	signal d_h2f_axi_master_rid                                             : std_logic_vector(11 downto 0);  -- mm_interconnect_0:d_h2f_axi_master_rid -> d:h2f_RID
	signal d_h2f_axi_master_rready                                          : std_logic;                      -- d:h2f_RREADY -> mm_interconnect_0:d_h2f_axi_master_rready
	signal d_h2f_axi_master_awlen                                           : std_logic_vector(3 downto 0);   -- d:h2f_AWLEN -> mm_interconnect_0:d_h2f_axi_master_awlen
	signal d_h2f_axi_master_wid                                             : std_logic_vector(11 downto 0);  -- d:h2f_WID -> mm_interconnect_0:d_h2f_axi_master_wid
	signal d_h2f_axi_master_arcache                                         : std_logic_vector(3 downto 0);   -- d:h2f_ARCACHE -> mm_interconnect_0:d_h2f_axi_master_arcache
	signal d_h2f_axi_master_wvalid                                          : std_logic;                      -- d:h2f_WVALID -> mm_interconnect_0:d_h2f_axi_master_wvalid
	signal d_h2f_axi_master_araddr                                          : std_logic_vector(29 downto 0);  -- d:h2f_ARADDR -> mm_interconnect_0:d_h2f_axi_master_araddr
	signal d_h2f_axi_master_arprot                                          : std_logic_vector(2 downto 0);   -- d:h2f_ARPROT -> mm_interconnect_0:d_h2f_axi_master_arprot
	signal d_h2f_axi_master_awprot                                          : std_logic_vector(2 downto 0);   -- d:h2f_AWPROT -> mm_interconnect_0:d_h2f_axi_master_awprot
	signal d_h2f_axi_master_wdata                                           : std_logic_vector(63 downto 0);  -- d:h2f_WDATA -> mm_interconnect_0:d_h2f_axi_master_wdata
	signal d_h2f_axi_master_arvalid                                         : std_logic;                      -- d:h2f_ARVALID -> mm_interconnect_0:d_h2f_axi_master_arvalid
	signal d_h2f_axi_master_awcache                                         : std_logic_vector(3 downto 0);   -- d:h2f_AWCACHE -> mm_interconnect_0:d_h2f_axi_master_awcache
	signal d_h2f_axi_master_arid                                            : std_logic_vector(11 downto 0);  -- d:h2f_ARID -> mm_interconnect_0:d_h2f_axi_master_arid
	signal d_h2f_axi_master_arlock                                          : std_logic_vector(1 downto 0);   -- d:h2f_ARLOCK -> mm_interconnect_0:d_h2f_axi_master_arlock
	signal d_h2f_axi_master_awlock                                          : std_logic_vector(1 downto 0);   -- d:h2f_AWLOCK -> mm_interconnect_0:d_h2f_axi_master_awlock
	signal d_h2f_axi_master_awaddr                                          : std_logic_vector(29 downto 0);  -- d:h2f_AWADDR -> mm_interconnect_0:d_h2f_axi_master_awaddr
	signal d_h2f_axi_master_bresp                                           : std_logic_vector(1 downto 0);   -- mm_interconnect_0:d_h2f_axi_master_bresp -> d:h2f_BRESP
	signal d_h2f_axi_master_arready                                         : std_logic;                      -- mm_interconnect_0:d_h2f_axi_master_arready -> d:h2f_ARREADY
	signal d_h2f_axi_master_rdata                                           : std_logic_vector(63 downto 0);  -- mm_interconnect_0:d_h2f_axi_master_rdata -> d:h2f_RDATA
	signal d_h2f_axi_master_awready                                         : std_logic;                      -- mm_interconnect_0:d_h2f_axi_master_awready -> d:h2f_AWREADY
	signal d_h2f_axi_master_arburst                                         : std_logic_vector(1 downto 0);   -- d:h2f_ARBURST -> mm_interconnect_0:d_h2f_axi_master_arburst
	signal d_h2f_axi_master_arsize                                          : std_logic_vector(2 downto 0);   -- d:h2f_ARSIZE -> mm_interconnect_0:d_h2f_axi_master_arsize
	signal d_h2f_axi_master_bready                                          : std_logic;                      -- d:h2f_BREADY -> mm_interconnect_0:d_h2f_axi_master_bready
	signal d_h2f_axi_master_rlast                                           : std_logic;                      -- mm_interconnect_0:d_h2f_axi_master_rlast -> d:h2f_RLAST
	signal d_h2f_axi_master_wlast                                           : std_logic;                      -- d:h2f_WLAST -> mm_interconnect_0:d_h2f_axi_master_wlast
	signal d_h2f_axi_master_rresp                                           : std_logic_vector(1 downto 0);   -- mm_interconnect_0:d_h2f_axi_master_rresp -> d:h2f_RRESP
	signal d_h2f_axi_master_awid                                            : std_logic_vector(11 downto 0);  -- d:h2f_AWID -> mm_interconnect_0:d_h2f_axi_master_awid
	signal d_h2f_axi_master_bid                                             : std_logic_vector(11 downto 0);  -- mm_interconnect_0:d_h2f_axi_master_bid -> d:h2f_BID
	signal d_h2f_axi_master_bvalid                                          : std_logic;                      -- mm_interconnect_0:d_h2f_axi_master_bvalid -> d:h2f_BVALID
	signal d_h2f_axi_master_awsize                                          : std_logic_vector(2 downto 0);   -- d:h2f_AWSIZE -> mm_interconnect_0:d_h2f_axi_master_awsize
	signal d_h2f_axi_master_awvalid                                         : std_logic;                      -- d:h2f_AWVALID -> mm_interconnect_0:d_h2f_axi_master_awvalid
	signal d_h2f_axi_master_rvalid                                          : std_logic;                      -- mm_interconnect_0:d_h2f_axi_master_rvalid -> d:h2f_RVALID
	signal fpga_only_master_master_readdata                                 : std_logic_vector(31 downto 0);  -- mm_interconnect_0:fpga_only_master_master_readdata -> fpga_only_master:master_readdata
	signal fpga_only_master_master_waitrequest                              : std_logic;                      -- mm_interconnect_0:fpga_only_master_master_waitrequest -> fpga_only_master:master_waitrequest
	signal fpga_only_master_master_address                                  : std_logic_vector(31 downto 0);  -- fpga_only_master:master_address -> mm_interconnect_0:fpga_only_master_master_address
	signal fpga_only_master_master_read                                     : std_logic;                      -- fpga_only_master:master_read -> mm_interconnect_0:fpga_only_master_master_read
	signal fpga_only_master_master_byteenable                               : std_logic_vector(3 downto 0);   -- fpga_only_master:master_byteenable -> mm_interconnect_0:fpga_only_master_master_byteenable
	signal fpga_only_master_master_readdatavalid                            : std_logic;                      -- mm_interconnect_0:fpga_only_master_master_readdatavalid -> fpga_only_master:master_readdatavalid
	signal fpga_only_master_master_write                                    : std_logic;                      -- fpga_only_master:master_write -> mm_interconnect_0:fpga_only_master_master_write
	signal fpga_only_master_master_writedata                                : std_logic_vector(31 downto 0);  -- fpga_only_master:master_writedata -> mm_interconnect_0:fpga_only_master_master_writedata
	signal d_h2f_lw_axi_master_awburst                                      : std_logic_vector(1 downto 0);   -- d:h2f_lw_AWBURST -> mm_interconnect_0:d_h2f_lw_axi_master_awburst
	signal d_h2f_lw_axi_master_arlen                                        : std_logic_vector(3 downto 0);   -- d:h2f_lw_ARLEN -> mm_interconnect_0:d_h2f_lw_axi_master_arlen
	signal d_h2f_lw_axi_master_wstrb                                        : std_logic_vector(3 downto 0);   -- d:h2f_lw_WSTRB -> mm_interconnect_0:d_h2f_lw_axi_master_wstrb
	signal d_h2f_lw_axi_master_wready                                       : std_logic;                      -- mm_interconnect_0:d_h2f_lw_axi_master_wready -> d:h2f_lw_WREADY
	signal d_h2f_lw_axi_master_rid                                          : std_logic_vector(11 downto 0);  -- mm_interconnect_0:d_h2f_lw_axi_master_rid -> d:h2f_lw_RID
	signal d_h2f_lw_axi_master_rready                                       : std_logic;                      -- d:h2f_lw_RREADY -> mm_interconnect_0:d_h2f_lw_axi_master_rready
	signal d_h2f_lw_axi_master_awlen                                        : std_logic_vector(3 downto 0);   -- d:h2f_lw_AWLEN -> mm_interconnect_0:d_h2f_lw_axi_master_awlen
	signal d_h2f_lw_axi_master_wid                                          : std_logic_vector(11 downto 0);  -- d:h2f_lw_WID -> mm_interconnect_0:d_h2f_lw_axi_master_wid
	signal d_h2f_lw_axi_master_arcache                                      : std_logic_vector(3 downto 0);   -- d:h2f_lw_ARCACHE -> mm_interconnect_0:d_h2f_lw_axi_master_arcache
	signal d_h2f_lw_axi_master_wvalid                                       : std_logic;                      -- d:h2f_lw_WVALID -> mm_interconnect_0:d_h2f_lw_axi_master_wvalid
	signal d_h2f_lw_axi_master_araddr                                       : std_logic_vector(20 downto 0);  -- d:h2f_lw_ARADDR -> mm_interconnect_0:d_h2f_lw_axi_master_araddr
	signal d_h2f_lw_axi_master_arprot                                       : std_logic_vector(2 downto 0);   -- d:h2f_lw_ARPROT -> mm_interconnect_0:d_h2f_lw_axi_master_arprot
	signal d_h2f_lw_axi_master_awprot                                       : std_logic_vector(2 downto 0);   -- d:h2f_lw_AWPROT -> mm_interconnect_0:d_h2f_lw_axi_master_awprot
	signal d_h2f_lw_axi_master_wdata                                        : std_logic_vector(31 downto 0);  -- d:h2f_lw_WDATA -> mm_interconnect_0:d_h2f_lw_axi_master_wdata
	signal d_h2f_lw_axi_master_arvalid                                      : std_logic;                      -- d:h2f_lw_ARVALID -> mm_interconnect_0:d_h2f_lw_axi_master_arvalid
	signal d_h2f_lw_axi_master_awcache                                      : std_logic_vector(3 downto 0);   -- d:h2f_lw_AWCACHE -> mm_interconnect_0:d_h2f_lw_axi_master_awcache
	signal d_h2f_lw_axi_master_arid                                         : std_logic_vector(11 downto 0);  -- d:h2f_lw_ARID -> mm_interconnect_0:d_h2f_lw_axi_master_arid
	signal d_h2f_lw_axi_master_arlock                                       : std_logic_vector(1 downto 0);   -- d:h2f_lw_ARLOCK -> mm_interconnect_0:d_h2f_lw_axi_master_arlock
	signal d_h2f_lw_axi_master_awlock                                       : std_logic_vector(1 downto 0);   -- d:h2f_lw_AWLOCK -> mm_interconnect_0:d_h2f_lw_axi_master_awlock
	signal d_h2f_lw_axi_master_awaddr                                       : std_logic_vector(20 downto 0);  -- d:h2f_lw_AWADDR -> mm_interconnect_0:d_h2f_lw_axi_master_awaddr
	signal d_h2f_lw_axi_master_bresp                                        : std_logic_vector(1 downto 0);   -- mm_interconnect_0:d_h2f_lw_axi_master_bresp -> d:h2f_lw_BRESP
	signal d_h2f_lw_axi_master_arready                                      : std_logic;                      -- mm_interconnect_0:d_h2f_lw_axi_master_arready -> d:h2f_lw_ARREADY
	signal d_h2f_lw_axi_master_rdata                                        : std_logic_vector(31 downto 0);  -- mm_interconnect_0:d_h2f_lw_axi_master_rdata -> d:h2f_lw_RDATA
	signal d_h2f_lw_axi_master_awready                                      : std_logic;                      -- mm_interconnect_0:d_h2f_lw_axi_master_awready -> d:h2f_lw_AWREADY
	signal d_h2f_lw_axi_master_arburst                                      : std_logic_vector(1 downto 0);   -- d:h2f_lw_ARBURST -> mm_interconnect_0:d_h2f_lw_axi_master_arburst
	signal d_h2f_lw_axi_master_arsize                                       : std_logic_vector(2 downto 0);   -- d:h2f_lw_ARSIZE -> mm_interconnect_0:d_h2f_lw_axi_master_arsize
	signal d_h2f_lw_axi_master_bready                                       : std_logic;                      -- d:h2f_lw_BREADY -> mm_interconnect_0:d_h2f_lw_axi_master_bready
	signal d_h2f_lw_axi_master_rlast                                        : std_logic;                      -- mm_interconnect_0:d_h2f_lw_axi_master_rlast -> d:h2f_lw_RLAST
	signal d_h2f_lw_axi_master_wlast                                        : std_logic;                      -- d:h2f_lw_WLAST -> mm_interconnect_0:d_h2f_lw_axi_master_wlast
	signal d_h2f_lw_axi_master_rresp                                        : std_logic_vector(1 downto 0);   -- mm_interconnect_0:d_h2f_lw_axi_master_rresp -> d:h2f_lw_RRESP
	signal d_h2f_lw_axi_master_awid                                         : std_logic_vector(11 downto 0);  -- d:h2f_lw_AWID -> mm_interconnect_0:d_h2f_lw_axi_master_awid
	signal d_h2f_lw_axi_master_bid                                          : std_logic_vector(11 downto 0);  -- mm_interconnect_0:d_h2f_lw_axi_master_bid -> d:h2f_lw_BID
	signal d_h2f_lw_axi_master_bvalid                                       : std_logic;                      -- mm_interconnect_0:d_h2f_lw_axi_master_bvalid -> d:h2f_lw_BVALID
	signal d_h2f_lw_axi_master_awsize                                       : std_logic_vector(2 downto 0);   -- d:h2f_lw_AWSIZE -> mm_interconnect_0:d_h2f_lw_axi_master_awsize
	signal d_h2f_lw_axi_master_awvalid                                      : std_logic;                      -- d:h2f_lw_AWVALID -> mm_interconnect_0:d_h2f_lw_axi_master_awvalid
	signal d_h2f_lw_axi_master_rvalid                                       : std_logic;                      -- mm_interconnect_0:d_h2f_lw_axi_master_rvalid -> d:h2f_lw_RVALID
	signal mm_interconnect_0_onchip_memory2_0_s1_chipselect                 : std_logic;                      -- mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	signal mm_interconnect_0_onchip_memory2_0_s1_readdata                   : std_logic_vector(63 downto 0);  -- onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	signal mm_interconnect_0_onchip_memory2_0_s1_address                    : std_logic_vector(12 downto 0);  -- mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	signal mm_interconnect_0_onchip_memory2_0_s1_byteenable                 : std_logic_vector(7 downto 0);   -- mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	signal mm_interconnect_0_onchip_memory2_0_s1_write                      : std_logic;                      -- mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	signal mm_interconnect_0_onchip_memory2_0_s1_writedata                  : std_logic_vector(63 downto 0);  -- mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_clken                      : std_logic;                      -- mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect         : std_logic;                      -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata           : std_logic_vector(31 downto 0);  -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest        : std_logic;                      -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address            : std_logic_vector(0 downto 0);   -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read               : std_logic;                      -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write              : std_logic;                      -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata          : std_logic_vector(31 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_intr_capturer_0_avalon_slave_0_readdata        : std_logic_vector(31 downto 0);  -- intr_capturer_0:rddata -> mm_interconnect_0:intr_capturer_0_avalon_slave_0_readdata
	signal mm_interconnect_0_intr_capturer_0_avalon_slave_0_address         : std_logic_vector(0 downto 0);   -- mm_interconnect_0:intr_capturer_0_avalon_slave_0_address -> intr_capturer_0:addr
	signal mm_interconnect_0_intr_capturer_0_avalon_slave_0_read            : std_logic;                      -- mm_interconnect_0:intr_capturer_0_avalon_slave_0_read -> intr_capturer_0:read
	signal mm_interconnect_0_sysid_qsys_control_slave_readdata              : std_logic_vector(31 downto 0);  -- sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	signal mm_interconnect_0_sysid_qsys_control_slave_address               : std_logic_vector(0 downto 0);   -- mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	signal mm_interconnect_0_led_pio_s1_chipselect                          : std_logic;                      -- mm_interconnect_0:led_pio_s1_chipselect -> led_pio:chipselect
	signal mm_interconnect_0_led_pio_s1_readdata                            : std_logic_vector(31 downto 0);  -- led_pio:readdata -> mm_interconnect_0:led_pio_s1_readdata
	signal mm_interconnect_0_led_pio_s1_address                             : std_logic_vector(1 downto 0);   -- mm_interconnect_0:led_pio_s1_address -> led_pio:address
	signal mm_interconnect_0_led_pio_s1_write                               : std_logic;                      -- mm_interconnect_0:led_pio_s1_write -> mm_interconnect_0_led_pio_s1_write:in
	signal mm_interconnect_0_led_pio_s1_writedata                           : std_logic_vector(31 downto 0);  -- mm_interconnect_0:led_pio_s1_writedata -> led_pio:writedata
	signal mm_interconnect_0_dipsw_pio_s1_chipselect                        : std_logic;                      -- mm_interconnect_0:dipsw_pio_s1_chipselect -> dipsw_pio:chipselect
	signal mm_interconnect_0_dipsw_pio_s1_readdata                          : std_logic_vector(31 downto 0);  -- dipsw_pio:readdata -> mm_interconnect_0:dipsw_pio_s1_readdata
	signal mm_interconnect_0_dipsw_pio_s1_address                           : std_logic_vector(1 downto 0);   -- mm_interconnect_0:dipsw_pio_s1_address -> dipsw_pio:address
	signal mm_interconnect_0_dipsw_pio_s1_write                             : std_logic;                      -- mm_interconnect_0:dipsw_pio_s1_write -> mm_interconnect_0_dipsw_pio_s1_write:in
	signal mm_interconnect_0_dipsw_pio_s1_writedata                         : std_logic_vector(31 downto 0);  -- mm_interconnect_0:dipsw_pio_s1_writedata -> dipsw_pio:writedata
	signal mm_interconnect_0_button_pio_s1_chipselect                       : std_logic;                      -- mm_interconnect_0:button_pio_s1_chipselect -> button_pio:chipselect
	signal mm_interconnect_0_button_pio_s1_readdata                         : std_logic_vector(31 downto 0);  -- button_pio:readdata -> mm_interconnect_0:button_pio_s1_readdata
	signal mm_interconnect_0_button_pio_s1_address                          : std_logic_vector(1 downto 0);   -- mm_interconnect_0:button_pio_s1_address -> button_pio:address
	signal mm_interconnect_0_button_pio_s1_write                            : std_logic;                      -- mm_interconnect_0:button_pio_s1_write -> mm_interconnect_0_button_pio_s1_write:in
	signal mm_interconnect_0_button_pio_s1_writedata                        : std_logic_vector(31 downto 0);  -- mm_interconnect_0:button_pio_s1_writedata -> button_pio:writedata
	signal mm_interconnect_0_ip_servomotor_0_avalon_slave_0_chipselect      : std_logic;                      -- mm_interconnect_0:IP_Servomotor_0_avalon_slave_0_chipselect -> IP_Servomotor_0:chip_select
	signal mm_interconnect_0_ip_servomotor_0_avalon_slave_0_address         : std_logic_vector(0 downto 0);   -- mm_interconnect_0:IP_Servomotor_0_avalon_slave_0_address -> IP_Servomotor_0:address
	signal mm_interconnect_0_ip_servomotor_0_avalon_slave_0_write           : std_logic;                      -- mm_interconnect_0:IP_Servomotor_0_avalon_slave_0_write -> mm_interconnect_0_ip_servomotor_0_avalon_slave_0_write:in
	signal mm_interconnect_0_ip_servomotor_0_avalon_slave_0_writedata       : std_logic_vector(7 downto 0);   -- mm_interconnect_0:IP_Servomotor_0_avalon_slave_0_writedata -> IP_Servomotor_0:write_data
	signal hps_only_master_master_readdata                                  : std_logic_vector(31 downto 0);  -- mm_interconnect_1:hps_only_master_master_readdata -> hps_only_master:master_readdata
	signal hps_only_master_master_waitrequest                               : std_logic;                      -- mm_interconnect_1:hps_only_master_master_waitrequest -> hps_only_master:master_waitrequest
	signal hps_only_master_master_address                                   : std_logic_vector(31 downto 0);  -- hps_only_master:master_address -> mm_interconnect_1:hps_only_master_master_address
	signal hps_only_master_master_read                                      : std_logic;                      -- hps_only_master:master_read -> mm_interconnect_1:hps_only_master_master_read
	signal hps_only_master_master_byteenable                                : std_logic_vector(3 downto 0);   -- hps_only_master:master_byteenable -> mm_interconnect_1:hps_only_master_master_byteenable
	signal hps_only_master_master_readdatavalid                             : std_logic;                      -- mm_interconnect_1:hps_only_master_master_readdatavalid -> hps_only_master:master_readdatavalid
	signal hps_only_master_master_write                                     : std_logic;                      -- hps_only_master:master_write -> mm_interconnect_1:hps_only_master_master_write
	signal hps_only_master_master_writedata                                 : std_logic_vector(31 downto 0);  -- hps_only_master:master_writedata -> mm_interconnect_1:hps_only_master_master_writedata
	signal mm_interconnect_1_d_f2h_axi_slave_awburst                        : std_logic_vector(1 downto 0);   -- mm_interconnect_1:d_f2h_axi_slave_awburst -> d:f2h_AWBURST
	signal mm_interconnect_1_d_f2h_axi_slave_awuser                         : std_logic_vector(4 downto 0);   -- mm_interconnect_1:d_f2h_axi_slave_awuser -> d:f2h_AWUSER
	signal mm_interconnect_1_d_f2h_axi_slave_arlen                          : std_logic_vector(3 downto 0);   -- mm_interconnect_1:d_f2h_axi_slave_arlen -> d:f2h_ARLEN
	signal mm_interconnect_1_d_f2h_axi_slave_wstrb                          : std_logic_vector(15 downto 0);  -- mm_interconnect_1:d_f2h_axi_slave_wstrb -> d:f2h_WSTRB
	signal mm_interconnect_1_d_f2h_axi_slave_wready                         : std_logic;                      -- d:f2h_WREADY -> mm_interconnect_1:d_f2h_axi_slave_wready
	signal mm_interconnect_1_d_f2h_axi_slave_rid                            : std_logic_vector(7 downto 0);   -- d:f2h_RID -> mm_interconnect_1:d_f2h_axi_slave_rid
	signal mm_interconnect_1_d_f2h_axi_slave_rready                         : std_logic;                      -- mm_interconnect_1:d_f2h_axi_slave_rready -> d:f2h_RREADY
	signal mm_interconnect_1_d_f2h_axi_slave_awlen                          : std_logic_vector(3 downto 0);   -- mm_interconnect_1:d_f2h_axi_slave_awlen -> d:f2h_AWLEN
	signal mm_interconnect_1_d_f2h_axi_slave_wid                            : std_logic_vector(7 downto 0);   -- mm_interconnect_1:d_f2h_axi_slave_wid -> d:f2h_WID
	signal mm_interconnect_1_d_f2h_axi_slave_arcache                        : std_logic_vector(3 downto 0);   -- mm_interconnect_1:d_f2h_axi_slave_arcache -> d:f2h_ARCACHE
	signal mm_interconnect_1_d_f2h_axi_slave_wvalid                         : std_logic;                      -- mm_interconnect_1:d_f2h_axi_slave_wvalid -> d:f2h_WVALID
	signal mm_interconnect_1_d_f2h_axi_slave_araddr                         : std_logic_vector(31 downto 0);  -- mm_interconnect_1:d_f2h_axi_slave_araddr -> d:f2h_ARADDR
	signal mm_interconnect_1_d_f2h_axi_slave_arprot                         : std_logic_vector(2 downto 0);   -- mm_interconnect_1:d_f2h_axi_slave_arprot -> d:f2h_ARPROT
	signal mm_interconnect_1_d_f2h_axi_slave_awprot                         : std_logic_vector(2 downto 0);   -- mm_interconnect_1:d_f2h_axi_slave_awprot -> d:f2h_AWPROT
	signal mm_interconnect_1_d_f2h_axi_slave_wdata                          : std_logic_vector(127 downto 0); -- mm_interconnect_1:d_f2h_axi_slave_wdata -> d:f2h_WDATA
	signal mm_interconnect_1_d_f2h_axi_slave_arvalid                        : std_logic;                      -- mm_interconnect_1:d_f2h_axi_slave_arvalid -> d:f2h_ARVALID
	signal mm_interconnect_1_d_f2h_axi_slave_awcache                        : std_logic_vector(3 downto 0);   -- mm_interconnect_1:d_f2h_axi_slave_awcache -> d:f2h_AWCACHE
	signal mm_interconnect_1_d_f2h_axi_slave_arid                           : std_logic_vector(7 downto 0);   -- mm_interconnect_1:d_f2h_axi_slave_arid -> d:f2h_ARID
	signal mm_interconnect_1_d_f2h_axi_slave_arlock                         : std_logic_vector(1 downto 0);   -- mm_interconnect_1:d_f2h_axi_slave_arlock -> d:f2h_ARLOCK
	signal mm_interconnect_1_d_f2h_axi_slave_awlock                         : std_logic_vector(1 downto 0);   -- mm_interconnect_1:d_f2h_axi_slave_awlock -> d:f2h_AWLOCK
	signal mm_interconnect_1_d_f2h_axi_slave_awaddr                         : std_logic_vector(31 downto 0);  -- mm_interconnect_1:d_f2h_axi_slave_awaddr -> d:f2h_AWADDR
	signal mm_interconnect_1_d_f2h_axi_slave_bresp                          : std_logic_vector(1 downto 0);   -- d:f2h_BRESP -> mm_interconnect_1:d_f2h_axi_slave_bresp
	signal mm_interconnect_1_d_f2h_axi_slave_arready                        : std_logic;                      -- d:f2h_ARREADY -> mm_interconnect_1:d_f2h_axi_slave_arready
	signal mm_interconnect_1_d_f2h_axi_slave_rdata                          : std_logic_vector(127 downto 0); -- d:f2h_RDATA -> mm_interconnect_1:d_f2h_axi_slave_rdata
	signal mm_interconnect_1_d_f2h_axi_slave_awready                        : std_logic;                      -- d:f2h_AWREADY -> mm_interconnect_1:d_f2h_axi_slave_awready
	signal mm_interconnect_1_d_f2h_axi_slave_arburst                        : std_logic_vector(1 downto 0);   -- mm_interconnect_1:d_f2h_axi_slave_arburst -> d:f2h_ARBURST
	signal mm_interconnect_1_d_f2h_axi_slave_arsize                         : std_logic_vector(2 downto 0);   -- mm_interconnect_1:d_f2h_axi_slave_arsize -> d:f2h_ARSIZE
	signal mm_interconnect_1_d_f2h_axi_slave_bready                         : std_logic;                      -- mm_interconnect_1:d_f2h_axi_slave_bready -> d:f2h_BREADY
	signal mm_interconnect_1_d_f2h_axi_slave_rlast                          : std_logic;                      -- d:f2h_RLAST -> mm_interconnect_1:d_f2h_axi_slave_rlast
	signal mm_interconnect_1_d_f2h_axi_slave_wlast                          : std_logic;                      -- mm_interconnect_1:d_f2h_axi_slave_wlast -> d:f2h_WLAST
	signal mm_interconnect_1_d_f2h_axi_slave_rresp                          : std_logic_vector(1 downto 0);   -- d:f2h_RRESP -> mm_interconnect_1:d_f2h_axi_slave_rresp
	signal mm_interconnect_1_d_f2h_axi_slave_awid                           : std_logic_vector(7 downto 0);   -- mm_interconnect_1:d_f2h_axi_slave_awid -> d:f2h_AWID
	signal mm_interconnect_1_d_f2h_axi_slave_bid                            : std_logic_vector(7 downto 0);   -- d:f2h_BID -> mm_interconnect_1:d_f2h_axi_slave_bid
	signal mm_interconnect_1_d_f2h_axi_slave_bvalid                         : std_logic;                      -- d:f2h_BVALID -> mm_interconnect_1:d_f2h_axi_slave_bvalid
	signal mm_interconnect_1_d_f2h_axi_slave_awsize                         : std_logic_vector(2 downto 0);   -- mm_interconnect_1:d_f2h_axi_slave_awsize -> d:f2h_AWSIZE
	signal mm_interconnect_1_d_f2h_axi_slave_awvalid                        : std_logic;                      -- mm_interconnect_1:d_f2h_axi_slave_awvalid -> d:f2h_AWVALID
	signal mm_interconnect_1_d_f2h_axi_slave_aruser                         : std_logic_vector(4 downto 0);   -- mm_interconnect_1:d_f2h_axi_slave_aruser -> d:f2h_ARUSER
	signal mm_interconnect_1_d_f2h_axi_slave_rvalid                         : std_logic;                      -- d:f2h_RVALID -> mm_interconnect_1:d_f2h_axi_slave_rvalid
	signal d_f2h_irq0_irq                                                   : std_logic_vector(31 downto 0);  -- irq_mapper:sender_irq -> d:f2h_irq_p0
	signal d_f2h_irq1_irq                                                   : std_logic_vector(31 downto 0);  -- irq_mapper_001:sender_irq -> d:f2h_irq_p1
	signal intr_capturer_0_interrupt_receiver_irq                           : std_logic_vector(31 downto 0);  -- irq_mapper_002:sender_irq -> intr_capturer_0:interrupt_in
	signal irq_mapper_receiver1_irq                                         : std_logic;                      -- button_pio:irq -> [irq_mapper:receiver1_irq, irq_mapper_002:receiver1_irq]
	signal irq_mapper_receiver2_irq                                         : std_logic;                      -- dipsw_pio:irq -> [irq_mapper:receiver2_irq, irq_mapper_002:receiver2_irq]
	signal irq_mapper_receiver0_irq                                         : std_logic;                      -- jtag_uart:av_irq -> [irq_mapper:receiver0_irq, irq_mapper_002:receiver0_irq]
	signal rst_controller_reset_out_reset                                   : std_logic;                      -- rst_controller:reset_out -> [irq_mapper_002:reset, mm_interconnect_0:fpga_only_master_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_0:onchip_memory2_0_reset1_reset_bridge_in_reset_reset, mm_interconnect_1:hps_only_master_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:hps_only_master_master_translator_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                               : std_logic;                      -- rst_controller:reset_req -> [onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	signal rst_controller_001_reset_out_reset                               : std_logic;                      -- rst_controller_001:reset_out -> [mm_interconnect_0:d_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:d_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset]
	signal hps_0_h2f_reset_reset_n_ports_inv                                : std_logic;                      -- hps_0_h2f_reset_reset_n:inv -> rst_controller_001:reset_in0
	signal reset_reset_n_ports_inv                                          : std_logic;                      -- reset_reset_n:inv -> [fpga_only_master:clk_reset_reset, hps_only_master:clk_reset_reset, rst_controller:reset_in0]
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv     : std_logic;                      -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv    : std_logic;                      -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_led_pio_s1_write_ports_inv                     : std_logic;                      -- mm_interconnect_0_led_pio_s1_write:inv -> led_pio:write_n
	signal mm_interconnect_0_dipsw_pio_s1_write_ports_inv                   : std_logic;                      -- mm_interconnect_0_dipsw_pio_s1_write:inv -> dipsw_pio:write_n
	signal mm_interconnect_0_button_pio_s1_write_ports_inv                  : std_logic;                      -- mm_interconnect_0_button_pio_s1_write:inv -> button_pio:write_n
	signal mm_interconnect_0_ip_servomotor_0_avalon_slave_0_write_ports_inv : std_logic;                      -- mm_interconnect_0_ip_servomotor_0_avalon_slave_0_write:inv -> IP_Servomotor_0:write_n
	signal rst_controller_reset_out_reset_ports_inv                         : std_logic;                      -- rst_controller_reset_out_reset:inv -> [IP_Servomotor_0:RST_n, button_pio:reset_n, dipsw_pio:reset_n, intr_capturer_0:rst_n, jtag_uart:rst_n, led_pio:reset_n, sysid_qsys:reset_n]

begin

	ip_servomotor_0 : component DF9GMS
		generic map (
			Fclock => 50000000
		)
		port map (
			address     => mm_interconnect_0_ip_servomotor_0_avalon_slave_0_address(0),      -- avalon_slave_0.address
			write_data  => mm_interconnect_0_ip_servomotor_0_avalon_slave_0_writedata,       --               .writedata
			write_n     => mm_interconnect_0_ip_servomotor_0_avalon_slave_0_write_ports_inv, --               .write_n
			chip_select => mm_interconnect_0_ip_servomotor_0_avalon_slave_0_chipselect,      --               .chipselect
			CLK         => clk_clk,                                                          --          clock.clk
			pulse       => ip_servomotor_0_conduit_end_commande,                             --    conduit_end.commande
			led         => ip_servomotor_0_conduit_end_led,                                  --               .led
			RST_n       => rst_controller_reset_out_reset_ports_inv                          --     reset_sink.reset_n
		);

	button_pio : component soc_system_button_pio
		port map (
			clk        => clk_clk,                                         --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,        --               reset.reset_n
			address    => mm_interconnect_0_button_pio_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_button_pio_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_button_pio_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_button_pio_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_button_pio_s1_readdata,        --                    .readdata
			in_port    => button_pio_external_connection_export,           -- external_connection.export
			irq        => irq_mapper_receiver1_irq                         --                 irq.irq
		);

	d : component soc_system_d
		generic map (
			F2S_Width => 3,
			S2F_Width => 2
		)
		port map (
			mem_a                    => memory_mem_a,                              --            memory.mem_a
			mem_ba                   => memory_mem_ba,                             --                  .mem_ba
			mem_ck                   => memory_mem_ck,                             --                  .mem_ck
			mem_ck_n                 => memory_mem_ck_n,                           --                  .mem_ck_n
			mem_cke                  => memory_mem_cke,                            --                  .mem_cke
			mem_cs_n                 => memory_mem_cs_n,                           --                  .mem_cs_n
			mem_ras_n                => memory_mem_ras_n,                          --                  .mem_ras_n
			mem_cas_n                => memory_mem_cas_n,                          --                  .mem_cas_n
			mem_we_n                 => memory_mem_we_n,                           --                  .mem_we_n
			mem_reset_n              => memory_mem_reset_n,                        --                  .mem_reset_n
			mem_dq                   => memory_mem_dq,                             --                  .mem_dq
			mem_dqs                  => memory_mem_dqs,                            --                  .mem_dqs
			mem_dqs_n                => memory_mem_dqs_n,                          --                  .mem_dqs_n
			mem_odt                  => memory_mem_odt,                            --                  .mem_odt
			mem_dm                   => memory_mem_dm,                             --                  .mem_dm
			oct_rzqin                => memory_oct_rzqin,                          --                  .oct_rzqin
			hps_io_emac1_inst_TX_CLK => hps_0_hps_io_hps_io_emac1_inst_TX_CLK,     --            hps_io.hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   => hps_0_hps_io_hps_io_emac1_inst_TXD0,       --                  .hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   => hps_0_hps_io_hps_io_emac1_inst_TXD1,       --                  .hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   => hps_0_hps_io_hps_io_emac1_inst_TXD2,       --                  .hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   => hps_0_hps_io_hps_io_emac1_inst_TXD3,       --                  .hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   => hps_0_hps_io_hps_io_emac1_inst_RXD0,       --                  .hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   => hps_0_hps_io_hps_io_emac1_inst_MDIO,       --                  .hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    => hps_0_hps_io_hps_io_emac1_inst_MDC,        --                  .hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL => hps_0_hps_io_hps_io_emac1_inst_RX_CTL,     --                  .hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL => hps_0_hps_io_hps_io_emac1_inst_TX_CTL,     --                  .hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK => hps_0_hps_io_hps_io_emac1_inst_RX_CLK,     --                  .hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   => hps_0_hps_io_hps_io_emac1_inst_RXD1,       --                  .hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   => hps_0_hps_io_hps_io_emac1_inst_RXD2,       --                  .hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   => hps_0_hps_io_hps_io_emac1_inst_RXD3,       --                  .hps_io_emac1_inst_RXD3
			hps_io_sdio_inst_CMD     => hps_0_hps_io_hps_io_sdio_inst_CMD,         --                  .hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      => hps_0_hps_io_hps_io_sdio_inst_D0,          --                  .hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      => hps_0_hps_io_hps_io_sdio_inst_D1,          --                  .hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     => hps_0_hps_io_hps_io_sdio_inst_CLK,         --                  .hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      => hps_0_hps_io_hps_io_sdio_inst_D2,          --                  .hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      => hps_0_hps_io_hps_io_sdio_inst_D3,          --                  .hps_io_sdio_inst_D3
			hps_io_usb1_inst_D0      => hps_0_hps_io_hps_io_usb1_inst_D0,          --                  .hps_io_usb1_inst_D0
			hps_io_usb1_inst_D1      => hps_0_hps_io_hps_io_usb1_inst_D1,          --                  .hps_io_usb1_inst_D1
			hps_io_usb1_inst_D2      => hps_0_hps_io_hps_io_usb1_inst_D2,          --                  .hps_io_usb1_inst_D2
			hps_io_usb1_inst_D3      => hps_0_hps_io_hps_io_usb1_inst_D3,          --                  .hps_io_usb1_inst_D3
			hps_io_usb1_inst_D4      => hps_0_hps_io_hps_io_usb1_inst_D4,          --                  .hps_io_usb1_inst_D4
			hps_io_usb1_inst_D5      => hps_0_hps_io_hps_io_usb1_inst_D5,          --                  .hps_io_usb1_inst_D5
			hps_io_usb1_inst_D6      => hps_0_hps_io_hps_io_usb1_inst_D6,          --                  .hps_io_usb1_inst_D6
			hps_io_usb1_inst_D7      => hps_0_hps_io_hps_io_usb1_inst_D7,          --                  .hps_io_usb1_inst_D7
			hps_io_usb1_inst_CLK     => hps_0_hps_io_hps_io_usb1_inst_CLK,         --                  .hps_io_usb1_inst_CLK
			hps_io_usb1_inst_STP     => hps_0_hps_io_hps_io_usb1_inst_STP,         --                  .hps_io_usb1_inst_STP
			hps_io_usb1_inst_DIR     => hps_0_hps_io_hps_io_usb1_inst_DIR,         --                  .hps_io_usb1_inst_DIR
			hps_io_usb1_inst_NXT     => hps_0_hps_io_hps_io_usb1_inst_NXT,         --                  .hps_io_usb1_inst_NXT
			hps_io_spim1_inst_CLK    => hps_0_hps_io_hps_io_spim1_inst_CLK,        --                  .hps_io_spim1_inst_CLK
			hps_io_spim1_inst_MOSI   => hps_0_hps_io_hps_io_spim1_inst_MOSI,       --                  .hps_io_spim1_inst_MOSI
			hps_io_spim1_inst_MISO   => hps_0_hps_io_hps_io_spim1_inst_MISO,       --                  .hps_io_spim1_inst_MISO
			hps_io_spim1_inst_SS0    => hps_0_hps_io_hps_io_spim1_inst_SS0,        --                  .hps_io_spim1_inst_SS0
			hps_io_uart0_inst_RX     => hps_0_hps_io_hps_io_uart0_inst_RX,         --                  .hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     => hps_0_hps_io_hps_io_uart0_inst_TX,         --                  .hps_io_uart0_inst_TX
			hps_io_i2c0_inst_SDA     => hps_0_hps_io_hps_io_i2c0_inst_SDA,         --                  .hps_io_i2c0_inst_SDA
			hps_io_i2c0_inst_SCL     => hps_0_hps_io_hps_io_i2c0_inst_SCL,         --                  .hps_io_i2c0_inst_SCL
			hps_io_i2c1_inst_SDA     => hps_0_hps_io_hps_io_i2c1_inst_SDA,         --                  .hps_io_i2c1_inst_SDA
			hps_io_i2c1_inst_SCL     => hps_0_hps_io_hps_io_i2c1_inst_SCL,         --                  .hps_io_i2c1_inst_SCL
			hps_io_gpio_inst_GPIO09  => hps_0_hps_io_hps_io_gpio_inst_GPIO09,      --                  .hps_io_gpio_inst_GPIO09
			hps_io_gpio_inst_GPIO35  => hps_0_hps_io_hps_io_gpio_inst_GPIO35,      --                  .hps_io_gpio_inst_GPIO35
			hps_io_gpio_inst_GPIO40  => hps_0_hps_io_hps_io_gpio_inst_GPIO40,      --                  .hps_io_gpio_inst_GPIO40
			hps_io_gpio_inst_GPIO53  => hps_0_hps_io_hps_io_gpio_inst_GPIO53,      --                  .hps_io_gpio_inst_GPIO53
			hps_io_gpio_inst_GPIO54  => hps_0_hps_io_hps_io_gpio_inst_GPIO54,      --                  .hps_io_gpio_inst_GPIO54
			hps_io_gpio_inst_GPIO61  => hps_0_hps_io_hps_io_gpio_inst_GPIO61,      --                  .hps_io_gpio_inst_GPIO61
			h2f_rst_n                => d_h2f_reset_reset,                         --         h2f_reset.reset_n
			h2f_axi_clk              => clk_clk,                                   --     h2f_axi_clock.clk
			h2f_AWID                 => d_h2f_axi_master_awid,                     --    h2f_axi_master.awid
			h2f_AWADDR               => d_h2f_axi_master_awaddr,                   --                  .awaddr
			h2f_AWLEN                => d_h2f_axi_master_awlen,                    --                  .awlen
			h2f_AWSIZE               => d_h2f_axi_master_awsize,                   --                  .awsize
			h2f_AWBURST              => d_h2f_axi_master_awburst,                  --                  .awburst
			h2f_AWLOCK               => d_h2f_axi_master_awlock,                   --                  .awlock
			h2f_AWCACHE              => d_h2f_axi_master_awcache,                  --                  .awcache
			h2f_AWPROT               => d_h2f_axi_master_awprot,                   --                  .awprot
			h2f_AWVALID              => d_h2f_axi_master_awvalid,                  --                  .awvalid
			h2f_AWREADY              => d_h2f_axi_master_awready,                  --                  .awready
			h2f_WID                  => d_h2f_axi_master_wid,                      --                  .wid
			h2f_WDATA                => d_h2f_axi_master_wdata,                    --                  .wdata
			h2f_WSTRB                => d_h2f_axi_master_wstrb,                    --                  .wstrb
			h2f_WLAST                => d_h2f_axi_master_wlast,                    --                  .wlast
			h2f_WVALID               => d_h2f_axi_master_wvalid,                   --                  .wvalid
			h2f_WREADY               => d_h2f_axi_master_wready,                   --                  .wready
			h2f_BID                  => d_h2f_axi_master_bid,                      --                  .bid
			h2f_BRESP                => d_h2f_axi_master_bresp,                    --                  .bresp
			h2f_BVALID               => d_h2f_axi_master_bvalid,                   --                  .bvalid
			h2f_BREADY               => d_h2f_axi_master_bready,                   --                  .bready
			h2f_ARID                 => d_h2f_axi_master_arid,                     --                  .arid
			h2f_ARADDR               => d_h2f_axi_master_araddr,                   --                  .araddr
			h2f_ARLEN                => d_h2f_axi_master_arlen,                    --                  .arlen
			h2f_ARSIZE               => d_h2f_axi_master_arsize,                   --                  .arsize
			h2f_ARBURST              => d_h2f_axi_master_arburst,                  --                  .arburst
			h2f_ARLOCK               => d_h2f_axi_master_arlock,                   --                  .arlock
			h2f_ARCACHE              => d_h2f_axi_master_arcache,                  --                  .arcache
			h2f_ARPROT               => d_h2f_axi_master_arprot,                   --                  .arprot
			h2f_ARVALID              => d_h2f_axi_master_arvalid,                  --                  .arvalid
			h2f_ARREADY              => d_h2f_axi_master_arready,                  --                  .arready
			h2f_RID                  => d_h2f_axi_master_rid,                      --                  .rid
			h2f_RDATA                => d_h2f_axi_master_rdata,                    --                  .rdata
			h2f_RRESP                => d_h2f_axi_master_rresp,                    --                  .rresp
			h2f_RLAST                => d_h2f_axi_master_rlast,                    --                  .rlast
			h2f_RVALID               => d_h2f_axi_master_rvalid,                   --                  .rvalid
			h2f_RREADY               => d_h2f_axi_master_rready,                   --                  .rready
			f2h_axi_clk              => clk_clk,                                   --     f2h_axi_clock.clk
			f2h_AWID                 => mm_interconnect_1_d_f2h_axi_slave_awid,    --     f2h_axi_slave.awid
			f2h_AWADDR               => mm_interconnect_1_d_f2h_axi_slave_awaddr,  --                  .awaddr
			f2h_AWLEN                => mm_interconnect_1_d_f2h_axi_slave_awlen,   --                  .awlen
			f2h_AWSIZE               => mm_interconnect_1_d_f2h_axi_slave_awsize,  --                  .awsize
			f2h_AWBURST              => mm_interconnect_1_d_f2h_axi_slave_awburst, --                  .awburst
			f2h_AWLOCK               => mm_interconnect_1_d_f2h_axi_slave_awlock,  --                  .awlock
			f2h_AWCACHE              => mm_interconnect_1_d_f2h_axi_slave_awcache, --                  .awcache
			f2h_AWPROT               => mm_interconnect_1_d_f2h_axi_slave_awprot,  --                  .awprot
			f2h_AWVALID              => mm_interconnect_1_d_f2h_axi_slave_awvalid, --                  .awvalid
			f2h_AWREADY              => mm_interconnect_1_d_f2h_axi_slave_awready, --                  .awready
			f2h_AWUSER               => mm_interconnect_1_d_f2h_axi_slave_awuser,  --                  .awuser
			f2h_WID                  => mm_interconnect_1_d_f2h_axi_slave_wid,     --                  .wid
			f2h_WDATA                => mm_interconnect_1_d_f2h_axi_slave_wdata,   --                  .wdata
			f2h_WSTRB                => mm_interconnect_1_d_f2h_axi_slave_wstrb,   --                  .wstrb
			f2h_WLAST                => mm_interconnect_1_d_f2h_axi_slave_wlast,   --                  .wlast
			f2h_WVALID               => mm_interconnect_1_d_f2h_axi_slave_wvalid,  --                  .wvalid
			f2h_WREADY               => mm_interconnect_1_d_f2h_axi_slave_wready,  --                  .wready
			f2h_BID                  => mm_interconnect_1_d_f2h_axi_slave_bid,     --                  .bid
			f2h_BRESP                => mm_interconnect_1_d_f2h_axi_slave_bresp,   --                  .bresp
			f2h_BVALID               => mm_interconnect_1_d_f2h_axi_slave_bvalid,  --                  .bvalid
			f2h_BREADY               => mm_interconnect_1_d_f2h_axi_slave_bready,  --                  .bready
			f2h_ARID                 => mm_interconnect_1_d_f2h_axi_slave_arid,    --                  .arid
			f2h_ARADDR               => mm_interconnect_1_d_f2h_axi_slave_araddr,  --                  .araddr
			f2h_ARLEN                => mm_interconnect_1_d_f2h_axi_slave_arlen,   --                  .arlen
			f2h_ARSIZE               => mm_interconnect_1_d_f2h_axi_slave_arsize,  --                  .arsize
			f2h_ARBURST              => mm_interconnect_1_d_f2h_axi_slave_arburst, --                  .arburst
			f2h_ARLOCK               => mm_interconnect_1_d_f2h_axi_slave_arlock,  --                  .arlock
			f2h_ARCACHE              => mm_interconnect_1_d_f2h_axi_slave_arcache, --                  .arcache
			f2h_ARPROT               => mm_interconnect_1_d_f2h_axi_slave_arprot,  --                  .arprot
			f2h_ARVALID              => mm_interconnect_1_d_f2h_axi_slave_arvalid, --                  .arvalid
			f2h_ARREADY              => mm_interconnect_1_d_f2h_axi_slave_arready, --                  .arready
			f2h_ARUSER               => mm_interconnect_1_d_f2h_axi_slave_aruser,  --                  .aruser
			f2h_RID                  => mm_interconnect_1_d_f2h_axi_slave_rid,     --                  .rid
			f2h_RDATA                => mm_interconnect_1_d_f2h_axi_slave_rdata,   --                  .rdata
			f2h_RRESP                => mm_interconnect_1_d_f2h_axi_slave_rresp,   --                  .rresp
			f2h_RLAST                => mm_interconnect_1_d_f2h_axi_slave_rlast,   --                  .rlast
			f2h_RVALID               => mm_interconnect_1_d_f2h_axi_slave_rvalid,  --                  .rvalid
			f2h_RREADY               => mm_interconnect_1_d_f2h_axi_slave_rready,  --                  .rready
			h2f_lw_axi_clk           => clk_clk,                                   --  h2f_lw_axi_clock.clk
			h2f_lw_AWID              => d_h2f_lw_axi_master_awid,                  -- h2f_lw_axi_master.awid
			h2f_lw_AWADDR            => d_h2f_lw_axi_master_awaddr,                --                  .awaddr
			h2f_lw_AWLEN             => d_h2f_lw_axi_master_awlen,                 --                  .awlen
			h2f_lw_AWSIZE            => d_h2f_lw_axi_master_awsize,                --                  .awsize
			h2f_lw_AWBURST           => d_h2f_lw_axi_master_awburst,               --                  .awburst
			h2f_lw_AWLOCK            => d_h2f_lw_axi_master_awlock,                --                  .awlock
			h2f_lw_AWCACHE           => d_h2f_lw_axi_master_awcache,               --                  .awcache
			h2f_lw_AWPROT            => d_h2f_lw_axi_master_awprot,                --                  .awprot
			h2f_lw_AWVALID           => d_h2f_lw_axi_master_awvalid,               --                  .awvalid
			h2f_lw_AWREADY           => d_h2f_lw_axi_master_awready,               --                  .awready
			h2f_lw_WID               => d_h2f_lw_axi_master_wid,                   --                  .wid
			h2f_lw_WDATA             => d_h2f_lw_axi_master_wdata,                 --                  .wdata
			h2f_lw_WSTRB             => d_h2f_lw_axi_master_wstrb,                 --                  .wstrb
			h2f_lw_WLAST             => d_h2f_lw_axi_master_wlast,                 --                  .wlast
			h2f_lw_WVALID            => d_h2f_lw_axi_master_wvalid,                --                  .wvalid
			h2f_lw_WREADY            => d_h2f_lw_axi_master_wready,                --                  .wready
			h2f_lw_BID               => d_h2f_lw_axi_master_bid,                   --                  .bid
			h2f_lw_BRESP             => d_h2f_lw_axi_master_bresp,                 --                  .bresp
			h2f_lw_BVALID            => d_h2f_lw_axi_master_bvalid,                --                  .bvalid
			h2f_lw_BREADY            => d_h2f_lw_axi_master_bready,                --                  .bready
			h2f_lw_ARID              => d_h2f_lw_axi_master_arid,                  --                  .arid
			h2f_lw_ARADDR            => d_h2f_lw_axi_master_araddr,                --                  .araddr
			h2f_lw_ARLEN             => d_h2f_lw_axi_master_arlen,                 --                  .arlen
			h2f_lw_ARSIZE            => d_h2f_lw_axi_master_arsize,                --                  .arsize
			h2f_lw_ARBURST           => d_h2f_lw_axi_master_arburst,               --                  .arburst
			h2f_lw_ARLOCK            => d_h2f_lw_axi_master_arlock,                --                  .arlock
			h2f_lw_ARCACHE           => d_h2f_lw_axi_master_arcache,               --                  .arcache
			h2f_lw_ARPROT            => d_h2f_lw_axi_master_arprot,                --                  .arprot
			h2f_lw_ARVALID           => d_h2f_lw_axi_master_arvalid,               --                  .arvalid
			h2f_lw_ARREADY           => d_h2f_lw_axi_master_arready,               --                  .arready
			h2f_lw_RID               => d_h2f_lw_axi_master_rid,                   --                  .rid
			h2f_lw_RDATA             => d_h2f_lw_axi_master_rdata,                 --                  .rdata
			h2f_lw_RRESP             => d_h2f_lw_axi_master_rresp,                 --                  .rresp
			h2f_lw_RLAST             => d_h2f_lw_axi_master_rlast,                 --                  .rlast
			h2f_lw_RVALID            => d_h2f_lw_axi_master_rvalid,                --                  .rvalid
			h2f_lw_RREADY            => d_h2f_lw_axi_master_rready,                --                  .rready
			f2h_irq_p0               => d_f2h_irq0_irq,                            --          f2h_irq0.irq
			f2h_irq_p1               => d_f2h_irq1_irq                             --          f2h_irq1.irq
		);

	dipsw_pio : component soc_system_dipsw_pio
		port map (
			clk        => clk_clk,                                        --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,       --               reset.reset_n
			address    => mm_interconnect_0_dipsw_pio_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_dipsw_pio_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_dipsw_pio_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_dipsw_pio_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_dipsw_pio_s1_readdata,        --                    .readdata
			in_port    => dipsw_pio_external_connection_export,           -- external_connection.export
			irq        => irq_mapper_receiver2_irq                        --                 irq.irq
		);

	fpga_only_master : component soc_system_fpga_only_master
		generic map (
			USE_PLI     => 0,
			PLI_PORT    => 50000,
			FIFO_DEPTHS => 2
		)
		port map (
			clk_clk              => clk_clk,                               --          clk.clk
			clk_reset_reset      => reset_reset_n_ports_inv,               --    clk_reset.reset
			master_address       => fpga_only_master_master_address,       --       master.address
			master_readdata      => fpga_only_master_master_readdata,      --             .readdata
			master_read          => fpga_only_master_master_read,          --             .read
			master_write         => fpga_only_master_master_write,         --             .write
			master_writedata     => fpga_only_master_master_writedata,     --             .writedata
			master_waitrequest   => fpga_only_master_master_waitrequest,   --             .waitrequest
			master_readdatavalid => fpga_only_master_master_readdatavalid, --             .readdatavalid
			master_byteenable    => fpga_only_master_master_byteenable,    --             .byteenable
			master_reset_reset   => open                                   -- master_reset.reset
		);

	hps_only_master : component soc_system_fpga_only_master
		generic map (
			USE_PLI     => 0,
			PLI_PORT    => 50000,
			FIFO_DEPTHS => 2
		)
		port map (
			clk_clk              => clk_clk,                              --          clk.clk
			clk_reset_reset      => reset_reset_n_ports_inv,              --    clk_reset.reset
			master_address       => hps_only_master_master_address,       --       master.address
			master_readdata      => hps_only_master_master_readdata,      --             .readdata
			master_read          => hps_only_master_master_read,          --             .read
			master_write         => hps_only_master_master_write,         --             .write
			master_writedata     => hps_only_master_master_writedata,     --             .writedata
			master_waitrequest   => hps_only_master_master_waitrequest,   --             .waitrequest
			master_readdatavalid => hps_only_master_master_readdatavalid, --             .readdatavalid
			master_byteenable    => hps_only_master_master_byteenable,    --             .byteenable
			master_reset_reset   => open                                  -- master_reset.reset
		);

	intr_capturer_0 : component intr_capturer
		generic map (
			NUM_INTR => 32
		)
		port map (
			clk          => clk_clk,                                                     --              clock.clk
			rst_n        => rst_controller_reset_out_reset_ports_inv,                    --         reset_sink.reset_n
			addr         => mm_interconnect_0_intr_capturer_0_avalon_slave_0_address(0), --     avalon_slave_0.address
			read         => mm_interconnect_0_intr_capturer_0_avalon_slave_0_read,       --                   .read
			rddata       => mm_interconnect_0_intr_capturer_0_avalon_slave_0_readdata,   --                   .readdata
			interrupt_in => intr_capturer_0_interrupt_receiver_irq                       -- interrupt_receiver.irq
		);

	jtag_uart : component soc_system_jtag_uart
		port map (
			clk            => clk_clk,                                                       --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                       --               irq.irq
		);

	led_pio : component soc_system_led_pio
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_led_pio_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_led_pio_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_led_pio_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_led_pio_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_led_pio_s1_readdata,        --                    .readdata
			out_port   => led_pio_external_connection_export            -- external_connection.export
		);

	onchip_memory2_0 : component soc_system_onchip_memory2_0
		port map (
			clk        => clk_clk,                                          --   clk1.clk
			address    => mm_interconnect_0_onchip_memory2_0_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory2_0_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory2_0_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory2_0_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory2_0_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory2_0_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory2_0_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                   -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,               --       .reset_req
			freeze     => '0'                                               -- (terminated)
		);

	sysid_qsys : component soc_system_sysid_qsys
		port map (
			clock    => clk_clk,                                               --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,              --         reset.reset_n
			readdata => mm_interconnect_0_sysid_qsys_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_qsys_control_slave_address(0)  --              .address
		);

	mm_interconnect_0 : component soc_system_mm_interconnect_0
		port map (
			d_h2f_axi_master_awid                                        => d_h2f_axi_master_awid,                                       --                                       d_h2f_axi_master.awid
			d_h2f_axi_master_awaddr                                      => d_h2f_axi_master_awaddr,                                     --                                                       .awaddr
			d_h2f_axi_master_awlen                                       => d_h2f_axi_master_awlen,                                      --                                                       .awlen
			d_h2f_axi_master_awsize                                      => d_h2f_axi_master_awsize,                                     --                                                       .awsize
			d_h2f_axi_master_awburst                                     => d_h2f_axi_master_awburst,                                    --                                                       .awburst
			d_h2f_axi_master_awlock                                      => d_h2f_axi_master_awlock,                                     --                                                       .awlock
			d_h2f_axi_master_awcache                                     => d_h2f_axi_master_awcache,                                    --                                                       .awcache
			d_h2f_axi_master_awprot                                      => d_h2f_axi_master_awprot,                                     --                                                       .awprot
			d_h2f_axi_master_awvalid                                     => d_h2f_axi_master_awvalid,                                    --                                                       .awvalid
			d_h2f_axi_master_awready                                     => d_h2f_axi_master_awready,                                    --                                                       .awready
			d_h2f_axi_master_wid                                         => d_h2f_axi_master_wid,                                        --                                                       .wid
			d_h2f_axi_master_wdata                                       => d_h2f_axi_master_wdata,                                      --                                                       .wdata
			d_h2f_axi_master_wstrb                                       => d_h2f_axi_master_wstrb,                                      --                                                       .wstrb
			d_h2f_axi_master_wlast                                       => d_h2f_axi_master_wlast,                                      --                                                       .wlast
			d_h2f_axi_master_wvalid                                      => d_h2f_axi_master_wvalid,                                     --                                                       .wvalid
			d_h2f_axi_master_wready                                      => d_h2f_axi_master_wready,                                     --                                                       .wready
			d_h2f_axi_master_bid                                         => d_h2f_axi_master_bid,                                        --                                                       .bid
			d_h2f_axi_master_bresp                                       => d_h2f_axi_master_bresp,                                      --                                                       .bresp
			d_h2f_axi_master_bvalid                                      => d_h2f_axi_master_bvalid,                                     --                                                       .bvalid
			d_h2f_axi_master_bready                                      => d_h2f_axi_master_bready,                                     --                                                       .bready
			d_h2f_axi_master_arid                                        => d_h2f_axi_master_arid,                                       --                                                       .arid
			d_h2f_axi_master_araddr                                      => d_h2f_axi_master_araddr,                                     --                                                       .araddr
			d_h2f_axi_master_arlen                                       => d_h2f_axi_master_arlen,                                      --                                                       .arlen
			d_h2f_axi_master_arsize                                      => d_h2f_axi_master_arsize,                                     --                                                       .arsize
			d_h2f_axi_master_arburst                                     => d_h2f_axi_master_arburst,                                    --                                                       .arburst
			d_h2f_axi_master_arlock                                      => d_h2f_axi_master_arlock,                                     --                                                       .arlock
			d_h2f_axi_master_arcache                                     => d_h2f_axi_master_arcache,                                    --                                                       .arcache
			d_h2f_axi_master_arprot                                      => d_h2f_axi_master_arprot,                                     --                                                       .arprot
			d_h2f_axi_master_arvalid                                     => d_h2f_axi_master_arvalid,                                    --                                                       .arvalid
			d_h2f_axi_master_arready                                     => d_h2f_axi_master_arready,                                    --                                                       .arready
			d_h2f_axi_master_rid                                         => d_h2f_axi_master_rid,                                        --                                                       .rid
			d_h2f_axi_master_rdata                                       => d_h2f_axi_master_rdata,                                      --                                                       .rdata
			d_h2f_axi_master_rresp                                       => d_h2f_axi_master_rresp,                                      --                                                       .rresp
			d_h2f_axi_master_rlast                                       => d_h2f_axi_master_rlast,                                      --                                                       .rlast
			d_h2f_axi_master_rvalid                                      => d_h2f_axi_master_rvalid,                                     --                                                       .rvalid
			d_h2f_axi_master_rready                                      => d_h2f_axi_master_rready,                                     --                                                       .rready
			d_h2f_lw_axi_master_awid                                     => d_h2f_lw_axi_master_awid,                                    --                                    d_h2f_lw_axi_master.awid
			d_h2f_lw_axi_master_awaddr                                   => d_h2f_lw_axi_master_awaddr,                                  --                                                       .awaddr
			d_h2f_lw_axi_master_awlen                                    => d_h2f_lw_axi_master_awlen,                                   --                                                       .awlen
			d_h2f_lw_axi_master_awsize                                   => d_h2f_lw_axi_master_awsize,                                  --                                                       .awsize
			d_h2f_lw_axi_master_awburst                                  => d_h2f_lw_axi_master_awburst,                                 --                                                       .awburst
			d_h2f_lw_axi_master_awlock                                   => d_h2f_lw_axi_master_awlock,                                  --                                                       .awlock
			d_h2f_lw_axi_master_awcache                                  => d_h2f_lw_axi_master_awcache,                                 --                                                       .awcache
			d_h2f_lw_axi_master_awprot                                   => d_h2f_lw_axi_master_awprot,                                  --                                                       .awprot
			d_h2f_lw_axi_master_awvalid                                  => d_h2f_lw_axi_master_awvalid,                                 --                                                       .awvalid
			d_h2f_lw_axi_master_awready                                  => d_h2f_lw_axi_master_awready,                                 --                                                       .awready
			d_h2f_lw_axi_master_wid                                      => d_h2f_lw_axi_master_wid,                                     --                                                       .wid
			d_h2f_lw_axi_master_wdata                                    => d_h2f_lw_axi_master_wdata,                                   --                                                       .wdata
			d_h2f_lw_axi_master_wstrb                                    => d_h2f_lw_axi_master_wstrb,                                   --                                                       .wstrb
			d_h2f_lw_axi_master_wlast                                    => d_h2f_lw_axi_master_wlast,                                   --                                                       .wlast
			d_h2f_lw_axi_master_wvalid                                   => d_h2f_lw_axi_master_wvalid,                                  --                                                       .wvalid
			d_h2f_lw_axi_master_wready                                   => d_h2f_lw_axi_master_wready,                                  --                                                       .wready
			d_h2f_lw_axi_master_bid                                      => d_h2f_lw_axi_master_bid,                                     --                                                       .bid
			d_h2f_lw_axi_master_bresp                                    => d_h2f_lw_axi_master_bresp,                                   --                                                       .bresp
			d_h2f_lw_axi_master_bvalid                                   => d_h2f_lw_axi_master_bvalid,                                  --                                                       .bvalid
			d_h2f_lw_axi_master_bready                                   => d_h2f_lw_axi_master_bready,                                  --                                                       .bready
			d_h2f_lw_axi_master_arid                                     => d_h2f_lw_axi_master_arid,                                    --                                                       .arid
			d_h2f_lw_axi_master_araddr                                   => d_h2f_lw_axi_master_araddr,                                  --                                                       .araddr
			d_h2f_lw_axi_master_arlen                                    => d_h2f_lw_axi_master_arlen,                                   --                                                       .arlen
			d_h2f_lw_axi_master_arsize                                   => d_h2f_lw_axi_master_arsize,                                  --                                                       .arsize
			d_h2f_lw_axi_master_arburst                                  => d_h2f_lw_axi_master_arburst,                                 --                                                       .arburst
			d_h2f_lw_axi_master_arlock                                   => d_h2f_lw_axi_master_arlock,                                  --                                                       .arlock
			d_h2f_lw_axi_master_arcache                                  => d_h2f_lw_axi_master_arcache,                                 --                                                       .arcache
			d_h2f_lw_axi_master_arprot                                   => d_h2f_lw_axi_master_arprot,                                  --                                                       .arprot
			d_h2f_lw_axi_master_arvalid                                  => d_h2f_lw_axi_master_arvalid,                                 --                                                       .arvalid
			d_h2f_lw_axi_master_arready                                  => d_h2f_lw_axi_master_arready,                                 --                                                       .arready
			d_h2f_lw_axi_master_rid                                      => d_h2f_lw_axi_master_rid,                                     --                                                       .rid
			d_h2f_lw_axi_master_rdata                                    => d_h2f_lw_axi_master_rdata,                                   --                                                       .rdata
			d_h2f_lw_axi_master_rresp                                    => d_h2f_lw_axi_master_rresp,                                   --                                                       .rresp
			d_h2f_lw_axi_master_rlast                                    => d_h2f_lw_axi_master_rlast,                                   --                                                       .rlast
			d_h2f_lw_axi_master_rvalid                                   => d_h2f_lw_axi_master_rvalid,                                  --                                                       .rvalid
			d_h2f_lw_axi_master_rready                                   => d_h2f_lw_axi_master_rready,                                  --                                                       .rready
			clk_0_clk_clk                                                => clk_clk,                                                     --                                              clk_0_clk.clk
			d_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                          -- d_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
			fpga_only_master_clk_reset_reset_bridge_in_reset_reset       => rst_controller_reset_out_reset,                              --       fpga_only_master_clk_reset_reset_bridge_in_reset.reset
			onchip_memory2_0_reset1_reset_bridge_in_reset_reset          => rst_controller_reset_out_reset,                              --          onchip_memory2_0_reset1_reset_bridge_in_reset.reset
			fpga_only_master_master_address                              => fpga_only_master_master_address,                             --                                fpga_only_master_master.address
			fpga_only_master_master_waitrequest                          => fpga_only_master_master_waitrequest,                         --                                                       .waitrequest
			fpga_only_master_master_byteenable                           => fpga_only_master_master_byteenable,                          --                                                       .byteenable
			fpga_only_master_master_read                                 => fpga_only_master_master_read,                                --                                                       .read
			fpga_only_master_master_readdata                             => fpga_only_master_master_readdata,                            --                                                       .readdata
			fpga_only_master_master_readdatavalid                        => fpga_only_master_master_readdatavalid,                       --                                                       .readdatavalid
			fpga_only_master_master_write                                => fpga_only_master_master_write,                               --                                                       .write
			fpga_only_master_master_writedata                            => fpga_only_master_master_writedata,                           --                                                       .writedata
			button_pio_s1_address                                        => mm_interconnect_0_button_pio_s1_address,                     --                                          button_pio_s1.address
			button_pio_s1_write                                          => mm_interconnect_0_button_pio_s1_write,                       --                                                       .write
			button_pio_s1_readdata                                       => mm_interconnect_0_button_pio_s1_readdata,                    --                                                       .readdata
			button_pio_s1_writedata                                      => mm_interconnect_0_button_pio_s1_writedata,                   --                                                       .writedata
			button_pio_s1_chipselect                                     => mm_interconnect_0_button_pio_s1_chipselect,                  --                                                       .chipselect
			dipsw_pio_s1_address                                         => mm_interconnect_0_dipsw_pio_s1_address,                      --                                           dipsw_pio_s1.address
			dipsw_pio_s1_write                                           => mm_interconnect_0_dipsw_pio_s1_write,                        --                                                       .write
			dipsw_pio_s1_readdata                                        => mm_interconnect_0_dipsw_pio_s1_readdata,                     --                                                       .readdata
			dipsw_pio_s1_writedata                                       => mm_interconnect_0_dipsw_pio_s1_writedata,                    --                                                       .writedata
			dipsw_pio_s1_chipselect                                      => mm_interconnect_0_dipsw_pio_s1_chipselect,                   --                                                       .chipselect
			intr_capturer_0_avalon_slave_0_address                       => mm_interconnect_0_intr_capturer_0_avalon_slave_0_address,    --                         intr_capturer_0_avalon_slave_0.address
			intr_capturer_0_avalon_slave_0_read                          => mm_interconnect_0_intr_capturer_0_avalon_slave_0_read,       --                                                       .read
			intr_capturer_0_avalon_slave_0_readdata                      => mm_interconnect_0_intr_capturer_0_avalon_slave_0_readdata,   --                                                       .readdata
			IP_Servomotor_0_avalon_slave_0_address                       => mm_interconnect_0_ip_servomotor_0_avalon_slave_0_address,    --                         IP_Servomotor_0_avalon_slave_0.address
			IP_Servomotor_0_avalon_slave_0_write                         => mm_interconnect_0_ip_servomotor_0_avalon_slave_0_write,      --                                                       .write
			IP_Servomotor_0_avalon_slave_0_writedata                     => mm_interconnect_0_ip_servomotor_0_avalon_slave_0_writedata,  --                                                       .writedata
			IP_Servomotor_0_avalon_slave_0_chipselect                    => mm_interconnect_0_ip_servomotor_0_avalon_slave_0_chipselect, --                                                       .chipselect
			jtag_uart_avalon_jtag_slave_address                          => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,       --                            jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write                            => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,         --                                                       .write
			jtag_uart_avalon_jtag_slave_read                             => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,          --                                                       .read
			jtag_uart_avalon_jtag_slave_readdata                         => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,      --                                                       .readdata
			jtag_uart_avalon_jtag_slave_writedata                        => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,     --                                                       .writedata
			jtag_uart_avalon_jtag_slave_waitrequest                      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,   --                                                       .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                       => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,    --                                                       .chipselect
			led_pio_s1_address                                           => mm_interconnect_0_led_pio_s1_address,                        --                                             led_pio_s1.address
			led_pio_s1_write                                             => mm_interconnect_0_led_pio_s1_write,                          --                                                       .write
			led_pio_s1_readdata                                          => mm_interconnect_0_led_pio_s1_readdata,                       --                                                       .readdata
			led_pio_s1_writedata                                         => mm_interconnect_0_led_pio_s1_writedata,                      --                                                       .writedata
			led_pio_s1_chipselect                                        => mm_interconnect_0_led_pio_s1_chipselect,                     --                                                       .chipselect
			onchip_memory2_0_s1_address                                  => mm_interconnect_0_onchip_memory2_0_s1_address,               --                                    onchip_memory2_0_s1.address
			onchip_memory2_0_s1_write                                    => mm_interconnect_0_onchip_memory2_0_s1_write,                 --                                                       .write
			onchip_memory2_0_s1_readdata                                 => mm_interconnect_0_onchip_memory2_0_s1_readdata,              --                                                       .readdata
			onchip_memory2_0_s1_writedata                                => mm_interconnect_0_onchip_memory2_0_s1_writedata,             --                                                       .writedata
			onchip_memory2_0_s1_byteenable                               => mm_interconnect_0_onchip_memory2_0_s1_byteenable,            --                                                       .byteenable
			onchip_memory2_0_s1_chipselect                               => mm_interconnect_0_onchip_memory2_0_s1_chipselect,            --                                                       .chipselect
			onchip_memory2_0_s1_clken                                    => mm_interconnect_0_onchip_memory2_0_s1_clken,                 --                                                       .clken
			sysid_qsys_control_slave_address                             => mm_interconnect_0_sysid_qsys_control_slave_address,          --                               sysid_qsys_control_slave.address
			sysid_qsys_control_slave_readdata                            => mm_interconnect_0_sysid_qsys_control_slave_readdata          --                                                       .readdata
		);

	mm_interconnect_1 : component soc_system_mm_interconnect_1
		port map (
			d_f2h_axi_slave_awid                                                => mm_interconnect_1_d_f2h_axi_slave_awid,    --                                               d_f2h_axi_slave.awid
			d_f2h_axi_slave_awaddr                                              => mm_interconnect_1_d_f2h_axi_slave_awaddr,  --                                                              .awaddr
			d_f2h_axi_slave_awlen                                               => mm_interconnect_1_d_f2h_axi_slave_awlen,   --                                                              .awlen
			d_f2h_axi_slave_awsize                                              => mm_interconnect_1_d_f2h_axi_slave_awsize,  --                                                              .awsize
			d_f2h_axi_slave_awburst                                             => mm_interconnect_1_d_f2h_axi_slave_awburst, --                                                              .awburst
			d_f2h_axi_slave_awlock                                              => mm_interconnect_1_d_f2h_axi_slave_awlock,  --                                                              .awlock
			d_f2h_axi_slave_awcache                                             => mm_interconnect_1_d_f2h_axi_slave_awcache, --                                                              .awcache
			d_f2h_axi_slave_awprot                                              => mm_interconnect_1_d_f2h_axi_slave_awprot,  --                                                              .awprot
			d_f2h_axi_slave_awuser                                              => mm_interconnect_1_d_f2h_axi_slave_awuser,  --                                                              .awuser
			d_f2h_axi_slave_awvalid                                             => mm_interconnect_1_d_f2h_axi_slave_awvalid, --                                                              .awvalid
			d_f2h_axi_slave_awready                                             => mm_interconnect_1_d_f2h_axi_slave_awready, --                                                              .awready
			d_f2h_axi_slave_wid                                                 => mm_interconnect_1_d_f2h_axi_slave_wid,     --                                                              .wid
			d_f2h_axi_slave_wdata                                               => mm_interconnect_1_d_f2h_axi_slave_wdata,   --                                                              .wdata
			d_f2h_axi_slave_wstrb                                               => mm_interconnect_1_d_f2h_axi_slave_wstrb,   --                                                              .wstrb
			d_f2h_axi_slave_wlast                                               => mm_interconnect_1_d_f2h_axi_slave_wlast,   --                                                              .wlast
			d_f2h_axi_slave_wvalid                                              => mm_interconnect_1_d_f2h_axi_slave_wvalid,  --                                                              .wvalid
			d_f2h_axi_slave_wready                                              => mm_interconnect_1_d_f2h_axi_slave_wready,  --                                                              .wready
			d_f2h_axi_slave_bid                                                 => mm_interconnect_1_d_f2h_axi_slave_bid,     --                                                              .bid
			d_f2h_axi_slave_bresp                                               => mm_interconnect_1_d_f2h_axi_slave_bresp,   --                                                              .bresp
			d_f2h_axi_slave_bvalid                                              => mm_interconnect_1_d_f2h_axi_slave_bvalid,  --                                                              .bvalid
			d_f2h_axi_slave_bready                                              => mm_interconnect_1_d_f2h_axi_slave_bready,  --                                                              .bready
			d_f2h_axi_slave_arid                                                => mm_interconnect_1_d_f2h_axi_slave_arid,    --                                                              .arid
			d_f2h_axi_slave_araddr                                              => mm_interconnect_1_d_f2h_axi_slave_araddr,  --                                                              .araddr
			d_f2h_axi_slave_arlen                                               => mm_interconnect_1_d_f2h_axi_slave_arlen,   --                                                              .arlen
			d_f2h_axi_slave_arsize                                              => mm_interconnect_1_d_f2h_axi_slave_arsize,  --                                                              .arsize
			d_f2h_axi_slave_arburst                                             => mm_interconnect_1_d_f2h_axi_slave_arburst, --                                                              .arburst
			d_f2h_axi_slave_arlock                                              => mm_interconnect_1_d_f2h_axi_slave_arlock,  --                                                              .arlock
			d_f2h_axi_slave_arcache                                             => mm_interconnect_1_d_f2h_axi_slave_arcache, --                                                              .arcache
			d_f2h_axi_slave_arprot                                              => mm_interconnect_1_d_f2h_axi_slave_arprot,  --                                                              .arprot
			d_f2h_axi_slave_aruser                                              => mm_interconnect_1_d_f2h_axi_slave_aruser,  --                                                              .aruser
			d_f2h_axi_slave_arvalid                                             => mm_interconnect_1_d_f2h_axi_slave_arvalid, --                                                              .arvalid
			d_f2h_axi_slave_arready                                             => mm_interconnect_1_d_f2h_axi_slave_arready, --                                                              .arready
			d_f2h_axi_slave_rid                                                 => mm_interconnect_1_d_f2h_axi_slave_rid,     --                                                              .rid
			d_f2h_axi_slave_rdata                                               => mm_interconnect_1_d_f2h_axi_slave_rdata,   --                                                              .rdata
			d_f2h_axi_slave_rresp                                               => mm_interconnect_1_d_f2h_axi_slave_rresp,   --                                                              .rresp
			d_f2h_axi_slave_rlast                                               => mm_interconnect_1_d_f2h_axi_slave_rlast,   --                                                              .rlast
			d_f2h_axi_slave_rvalid                                              => mm_interconnect_1_d_f2h_axi_slave_rvalid,  --                                                              .rvalid
			d_f2h_axi_slave_rready                                              => mm_interconnect_1_d_f2h_axi_slave_rready,  --                                                              .rready
			clk_0_clk_clk                                                       => clk_clk,                                   --                                                     clk_0_clk.clk
			d_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset        => rst_controller_001_reset_out_reset,        --        d_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset.reset
			hps_only_master_clk_reset_reset_bridge_in_reset_reset               => rst_controller_reset_out_reset,            --               hps_only_master_clk_reset_reset_bridge_in_reset.reset
			hps_only_master_master_translator_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,            -- hps_only_master_master_translator_reset_reset_bridge_in_reset.reset
			hps_only_master_master_address                                      => hps_only_master_master_address,            --                                        hps_only_master_master.address
			hps_only_master_master_waitrequest                                  => hps_only_master_master_waitrequest,        --                                                              .waitrequest
			hps_only_master_master_byteenable                                   => hps_only_master_master_byteenable,         --                                                              .byteenable
			hps_only_master_master_read                                         => hps_only_master_master_read,               --                                                              .read
			hps_only_master_master_readdata                                     => hps_only_master_master_readdata,           --                                                              .readdata
			hps_only_master_master_readdatavalid                                => hps_only_master_master_readdatavalid,      --                                                              .readdatavalid
			hps_only_master_master_write                                        => hps_only_master_master_write,              --                                                              .write
			hps_only_master_master_writedata                                    => hps_only_master_master_writedata           --                                                              .writedata
		);

	irq_mapper : component soc_system_irq_mapper
		port map (
			clk           => open,                     --       clk.clk
			reset         => open,                     -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq, -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq, -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq, -- receiver2.irq
			sender_irq    => d_f2h_irq0_irq            --    sender.irq
		);

	irq_mapper_001 : component soc_system_irq_mapper_001
		port map (
			clk        => open,           --       clk.clk
			reset      => open,           -- clk_reset.reset
			sender_irq => d_f2h_irq1_irq  --    sender.irq
		);

	irq_mapper_002 : component soc_system_irq_mapper
		port map (
			clk           => clk_clk,                                --       clk.clk
			reset         => rst_controller_reset_out_reset,         -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,               -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,               -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,               -- receiver2.irq
			sender_irq    => intr_capturer_0_interrupt_receiver_irq  --    sender.irq
		);

	rst_controller : component soc_system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component soc_system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => hps_0_h2f_reset_reset_n_ports_inv,  -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	hps_0_h2f_reset_reset_n_ports_inv <= not d_h2f_reset_reset;

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_led_pio_s1_write_ports_inv <= not mm_interconnect_0_led_pio_s1_write;

	mm_interconnect_0_dipsw_pio_s1_write_ports_inv <= not mm_interconnect_0_dipsw_pio_s1_write;

	mm_interconnect_0_button_pio_s1_write_ports_inv <= not mm_interconnect_0_button_pio_s1_write;

	mm_interconnect_0_ip_servomotor_0_avalon_slave_0_write_ports_inv <= not mm_interconnect_0_ip_servomotor_0_avalon_slave_0_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	hps_0_h2f_reset_reset_n <= d_h2f_reset_reset;

end architecture rtl; -- of soc_system
